// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : mul_4
// Git hash  : fbf001df014e844f818dd31ebd5c3686888b43b3


module mul_4 (
  input      [63:0]   A,
  input      [63:0]   B,
  output     [63:0]   P,
  input               clk,
  input               reset
);
  wire       [127:0]  _zz_P_6;
  (* use_dsp = "yes" *) wire       [63:0]   _zz_P;
  (* use_dsp = "yes" *) wire       [63:0]   _zz_P_1;
  (* use_dsp = "yes" *) reg        [63:0]   _zz_P_2;
  (* use_dsp = "yes" *) reg        [63:0]   _zz_P_3;
  (* use_dsp = "yes" *) reg        [127:0]  _zz_P_4;
  (* use_dsp = "yes" *) reg        [127:0]  _zz_P_5;

  assign _zz_P_6 = _zz_P_5;
  assign _zz_P = A;
  assign _zz_P_1 = B;
  assign P = _zz_P_6[63:0];
  always @(posedge clk) begin
    _zz_P_2 <= _zz_P;
    _zz_P_3 <= _zz_P_1;
    _zz_P_4 <= (_zz_P_2 * _zz_P_3);
    _zz_P_5 <= _zz_P_4;
  end


endmodule
