// Generator : SpinalHDL v1.4.3    git head : adf552d8f500e7419fff395b7049228e4bc5de26
// Component : TestEnv
// Git hash  : 6b765f9792de40c223ec28811737ae22b58a9fa8



module TestEnv (
  input               a,
  output              b
);

  assign b = a;

endmodule
