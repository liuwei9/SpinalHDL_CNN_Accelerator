// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : A
// Git hash  : b694a57c8f5c199d7fd0af5809d5f7d2954eb351



module A (
  input               _zz_1,
  output              _zz_2
);

  assign _zz_2 = _zz_1;

endmodule
