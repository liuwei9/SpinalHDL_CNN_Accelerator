// Generator : SpinalHDL v1.6.0    git head : 73c8d8e2b86b45646e9d0b2e729291f2b65e6be3
// Component : Conv_Norm
// Git hash  : a7a69259854496944a80b53cb839562d830e2b39
// Date      : 17/09/2021, 17:43:46


module Conv_Norm (
  input               Start_Cu,
  input               Start_Pa,
  input               para_data_valid,
  output              para_data_ready,
  input      [63:0]   para_data_payload,
  output              Write_Block_Complete,
  output              Compute_Complete,
  input      [575:0]  S_DATA,
  input      [8:0]    S_DATA_Valid,
  output              S_DATA_Ready,
  output reg          M_DATA_valid,
  input               M_DATA_ready,
  output reg [255:0]  M_DATA_payload,
  input      [10:0]   Row_Num_Out_REG,
  input      [10:0]   RowNum_After_Padding,
  input      [9:0]    Channel_In_Num_REG,
  input      [9:0]    Channel_Out_Num_REG,
  input      [14:0]   Weight_Single_Num_REG,
  input      [7:0]    Bias_Num_REG,
  input      [7:0]    Bias_Addrb,
  output     [255:0]  Data_Out_Bias,
  output     [255:0]  Data_Out_Scale,
  output     [255:0]  Data_Out_Shift,
  input               clk,
  input               reset
);
  wire                compute_ctrl_1_compute_fifo_ready;
  wire       [10:0]   compute_ctrl_1_COMPUTE_TIMES_CHANNEL_IN_REG;
  wire       [10:0]   compute_ctrl_1_COMPUTE_TIMES_CHANNEL_IN_REG_8;
  wire       [10:0]   compute_ctrl_1_COMPUTE_TIMES_CHANNEL_OUT_REG;
  wire       [63:0]   general_fifo_sync_10_data_in;
  wire                general_fifo_sync_10_wr_en;
  wire       [10:0]   general_fifo_sync_10_m_data_count;
  wire       [10:0]   general_fifo_sync_10_s_data_count;
  wire       [63:0]   general_fifo_sync_11_data_in;
  wire                general_fifo_sync_11_wr_en;
  wire       [10:0]   general_fifo_sync_11_m_data_count;
  wire       [10:0]   general_fifo_sync_11_s_data_count;
  wire       [63:0]   general_fifo_sync_12_data_in;
  wire                general_fifo_sync_12_wr_en;
  wire       [10:0]   general_fifo_sync_12_m_data_count;
  wire       [10:0]   general_fifo_sync_12_s_data_count;
  wire       [63:0]   general_fifo_sync_13_data_in;
  wire                general_fifo_sync_13_wr_en;
  wire       [10:0]   general_fifo_sync_13_m_data_count;
  wire       [10:0]   general_fifo_sync_13_s_data_count;
  wire       [63:0]   general_fifo_sync_14_data_in;
  wire                general_fifo_sync_14_wr_en;
  wire       [10:0]   general_fifo_sync_14_m_data_count;
  wire       [10:0]   general_fifo_sync_14_s_data_count;
  wire       [63:0]   general_fifo_sync_15_data_in;
  wire                general_fifo_sync_15_wr_en;
  wire       [10:0]   general_fifo_sync_15_m_data_count;
  wire       [10:0]   general_fifo_sync_15_s_data_count;
  wire       [63:0]   general_fifo_sync_16_data_in;
  wire                general_fifo_sync_16_wr_en;
  wire       [10:0]   general_fifo_sync_16_m_data_count;
  wire       [10:0]   general_fifo_sync_16_s_data_count;
  wire       [63:0]   general_fifo_sync_17_data_in;
  wire                general_fifo_sync_17_wr_en;
  wire       [10:0]   general_fifo_sync_17_m_data_count;
  wire       [10:0]   general_fifo_sync_17_s_data_count;
  wire       [63:0]   general_fifo_sync_18_data_in;
  wire                general_fifo_sync_18_wr_en;
  wire       [10:0]   general_fifo_sync_18_m_data_count;
  wire       [10:0]   general_fifo_sync_18_s_data_count;
  wire       [0:0]    Configurable_RAM_Norm_wea;
  wire       [71:0]   mul_add_simd_128_weightIn;
  wire       [71:0]   mul_add_simd_129_weightIn;
  wire       [71:0]   mul_add_simd_130_weightIn;
  wire       [71:0]   mul_add_simd_131_weightIn;
  wire       [71:0]   mul_add_simd_132_weightIn;
  wire       [71:0]   mul_add_simd_133_weightIn;
  wire       [71:0]   mul_add_simd_134_weightIn;
  wire       [71:0]   mul_add_simd_135_weightIn;
  wire       [71:0]   mul_add_simd_136_weightIn;
  wire       [71:0]   mul_add_simd_137_weightIn;
  wire       [71:0]   mul_add_simd_138_weightIn;
  wire       [71:0]   mul_add_simd_139_weightIn;
  wire       [71:0]   mul_add_simd_140_weightIn;
  wire       [71:0]   mul_add_simd_141_weightIn;
  wire       [71:0]   mul_add_simd_142_weightIn;
  wire       [71:0]   mul_add_simd_143_weightIn;
  wire       [71:0]   mul_add_simd_144_weightIn;
  wire       [71:0]   mul_add_simd_145_weightIn;
  wire       [71:0]   mul_add_simd_146_weightIn;
  wire       [71:0]   mul_add_simd_147_weightIn;
  wire       [71:0]   mul_add_simd_148_weightIn;
  wire       [71:0]   mul_add_simd_149_weightIn;
  wire       [71:0]   mul_add_simd_150_weightIn;
  wire       [71:0]   mul_add_simd_151_weightIn;
  wire       [71:0]   mul_add_simd_152_weightIn;
  wire       [71:0]   mul_add_simd_153_weightIn;
  wire       [71:0]   mul_add_simd_154_weightIn;
  wire       [71:0]   mul_add_simd_155_weightIn;
  wire       [71:0]   mul_add_simd_156_weightIn;
  wire       [71:0]   mul_add_simd_157_weightIn;
  wire       [71:0]   mul_add_simd_158_weightIn;
  wire       [71:0]   mul_add_simd_159_weightIn;
  wire       [71:0]   mul_add_simd_160_weightIn;
  wire       [71:0]   mul_add_simd_161_weightIn;
  wire       [71:0]   mul_add_simd_162_weightIn;
  wire       [71:0]   mul_add_simd_163_weightIn;
  wire       [71:0]   mul_add_simd_164_weightIn;
  wire       [71:0]   mul_add_simd_165_weightIn;
  wire       [71:0]   mul_add_simd_166_weightIn;
  wire       [71:0]   mul_add_simd_167_weightIn;
  wire       [71:0]   mul_add_simd_168_weightIn;
  wire       [71:0]   mul_add_simd_169_weightIn;
  wire       [71:0]   mul_add_simd_170_weightIn;
  wire       [71:0]   mul_add_simd_171_weightIn;
  wire       [71:0]   mul_add_simd_172_weightIn;
  wire       [71:0]   mul_add_simd_173_weightIn;
  wire       [71:0]   mul_add_simd_174_weightIn;
  wire       [71:0]   mul_add_simd_175_weightIn;
  wire       [71:0]   mul_add_simd_176_weightIn;
  wire       [71:0]   mul_add_simd_177_weightIn;
  wire       [71:0]   mul_add_simd_178_weightIn;
  wire       [71:0]   mul_add_simd_179_weightIn;
  wire       [71:0]   mul_add_simd_180_weightIn;
  wire       [71:0]   mul_add_simd_181_weightIn;
  wire       [71:0]   mul_add_simd_182_weightIn;
  wire       [71:0]   mul_add_simd_183_weightIn;
  wire       [71:0]   mul_add_simd_184_weightIn;
  wire       [71:0]   mul_add_simd_185_weightIn;
  wire       [71:0]   mul_add_simd_186_weightIn;
  wire       [71:0]   mul_add_simd_187_weightIn;
  wire       [71:0]   mul_add_simd_188_weightIn;
  wire       [71:0]   mul_add_simd_189_weightIn;
  wire       [71:0]   mul_add_simd_190_weightIn;
  wire       [71:0]   mul_add_simd_191_weightIn;
  wire       [71:0]   mul_add_simd_192_weightIn;
  wire       [71:0]   mul_add_simd_193_weightIn;
  wire       [71:0]   mul_add_simd_194_weightIn;
  wire       [71:0]   mul_add_simd_195_weightIn;
  wire       [71:0]   mul_add_simd_196_weightIn;
  wire       [71:0]   mul_add_simd_197_weightIn;
  wire       [71:0]   mul_add_simd_198_weightIn;
  wire       [71:0]   mul_add_simd_199_weightIn;
  wire       [71:0]   mul_add_simd_200_weightIn;
  wire       [71:0]   mul_add_simd_201_weightIn;
  wire       [71:0]   mul_add_simd_202_weightIn;
  wire       [71:0]   mul_add_simd_203_weightIn;
  wire       [71:0]   mul_add_simd_204_weightIn;
  wire       [71:0]   mul_add_simd_205_weightIn;
  wire       [71:0]   mul_add_simd_206_weightIn;
  wire       [71:0]   mul_add_simd_207_weightIn;
  wire       [71:0]   mul_add_simd_208_weightIn;
  wire       [71:0]   mul_add_simd_209_weightIn;
  wire       [71:0]   mul_add_simd_210_weightIn;
  wire       [71:0]   mul_add_simd_211_weightIn;
  wire       [71:0]   mul_add_simd_212_weightIn;
  wire       [71:0]   mul_add_simd_213_weightIn;
  wire       [71:0]   mul_add_simd_214_weightIn;
  wire       [71:0]   mul_add_simd_215_weightIn;
  wire       [71:0]   mul_add_simd_216_weightIn;
  wire       [71:0]   mul_add_simd_217_weightIn;
  wire       [71:0]   mul_add_simd_218_weightIn;
  wire       [71:0]   mul_add_simd_219_weightIn;
  wire       [71:0]   mul_add_simd_220_weightIn;
  wire       [71:0]   mul_add_simd_221_weightIn;
  wire       [71:0]   mul_add_simd_222_weightIn;
  wire       [71:0]   mul_add_simd_223_weightIn;
  wire       [71:0]   mul_add_simd_224_weightIn;
  wire       [71:0]   mul_add_simd_225_weightIn;
  wire       [71:0]   mul_add_simd_226_weightIn;
  wire       [71:0]   mul_add_simd_227_weightIn;
  wire       [71:0]   mul_add_simd_228_weightIn;
  wire       [71:0]   mul_add_simd_229_weightIn;
  wire       [71:0]   mul_add_simd_230_weightIn;
  wire       [71:0]   mul_add_simd_231_weightIn;
  wire       [71:0]   mul_add_simd_232_weightIn;
  wire       [71:0]   mul_add_simd_233_weightIn;
  wire       [71:0]   mul_add_simd_234_weightIn;
  wire       [71:0]   mul_add_simd_235_weightIn;
  wire       [71:0]   mul_add_simd_236_weightIn;
  wire       [71:0]   mul_add_simd_237_weightIn;
  wire       [71:0]   mul_add_simd_238_weightIn;
  wire       [71:0]   mul_add_simd_239_weightIn;
  wire       [71:0]   mul_add_simd_240_weightIn;
  wire       [71:0]   mul_add_simd_241_weightIn;
  wire       [71:0]   mul_add_simd_242_weightIn;
  wire       [71:0]   mul_add_simd_243_weightIn;
  wire       [71:0]   mul_add_simd_244_weightIn;
  wire       [71:0]   mul_add_simd_245_weightIn;
  wire       [71:0]   mul_add_simd_246_weightIn;
  wire       [71:0]   mul_add_simd_247_weightIn;
  wire       [71:0]   mul_add_simd_248_weightIn;
  wire       [71:0]   mul_add_simd_249_weightIn;
  wire       [71:0]   mul_add_simd_250_weightIn;
  wire       [71:0]   mul_add_simd_251_weightIn;
  wire       [71:0]   mul_add_simd_252_weightIn;
  wire       [71:0]   mul_add_simd_253_weightIn;
  wire       [71:0]   mul_add_simd_254_weightIn;
  wire       [71:0]   mul_add_simd_255_weightIn;
  wire                compute_ctrl_1_Compute_Complete;
  wire                compute_ctrl_1_First_Compute_Complete;
  wire                compute_ctrl_1_rd_en_fifo;
  wire                compute_ctrl_1_M_Valid;
  wire       [12:0]   compute_ctrl_1_weight_addrb;
  wire       [10:0]   compute_ctrl_1_ram_temp_read_address;
  wire       [10:0]   compute_ctrl_1_ram_temp_write_address;
  wire       [10:0]   compute_ctrl_1_S_Count_Fifo;
  wire       [10:0]   compute_ctrl_1_M_Count_Fifo;
  wire                load_weight_1_Write_Block_Complete;
  wire                load_weight_1_S_Para_Data_ready;
  wire       [1023:0] load_weight_1_Data_Out_Weight_0;
  wire       [1023:0] load_weight_1_Data_Out_Weight_1;
  wire       [1023:0] load_weight_1_Data_Out_Weight_2;
  wire       [1023:0] load_weight_1_Data_Out_Weight_3;
  wire       [1023:0] load_weight_1_Data_Out_Weight_4;
  wire       [1023:0] load_weight_1_Data_Out_Weight_5;
  wire       [1023:0] load_weight_1_Data_Out_Weight_6;
  wire       [1023:0] load_weight_1_Data_Out_Weight_7;
  wire       [1023:0] load_weight_1_Data_Out_Weight_8;
  wire       [255:0]  load_weight_1_Data_Out_Bias;
  wire       [255:0]  load_weight_1_Data_Out_Scale;
  wire       [255:0]  load_weight_1_Data_Out_Shift;
  wire                general_fifo_sync_10_data_in_ready;
  wire       [127:0]  general_fifo_sync_10_data_out;
  wire                general_fifo_sync_10_data_out_valid;
  wire                general_fifo_sync_10_data_valid;
  wire                general_fifo_sync_10_full;
  wire                general_fifo_sync_10_empty;
  wire                general_fifo_sync_11_data_in_ready;
  wire       [127:0]  general_fifo_sync_11_data_out;
  wire                general_fifo_sync_11_data_out_valid;
  wire                general_fifo_sync_11_data_valid;
  wire                general_fifo_sync_11_full;
  wire                general_fifo_sync_11_empty;
  wire                general_fifo_sync_12_data_in_ready;
  wire       [127:0]  general_fifo_sync_12_data_out;
  wire                general_fifo_sync_12_data_out_valid;
  wire                general_fifo_sync_12_data_valid;
  wire                general_fifo_sync_12_full;
  wire                general_fifo_sync_12_empty;
  wire                general_fifo_sync_13_data_in_ready;
  wire       [127:0]  general_fifo_sync_13_data_out;
  wire                general_fifo_sync_13_data_out_valid;
  wire                general_fifo_sync_13_data_valid;
  wire                general_fifo_sync_13_full;
  wire                general_fifo_sync_13_empty;
  wire                general_fifo_sync_14_data_in_ready;
  wire       [127:0]  general_fifo_sync_14_data_out;
  wire                general_fifo_sync_14_data_out_valid;
  wire                general_fifo_sync_14_data_valid;
  wire                general_fifo_sync_14_full;
  wire                general_fifo_sync_14_empty;
  wire                general_fifo_sync_15_data_in_ready;
  wire       [127:0]  general_fifo_sync_15_data_out;
  wire                general_fifo_sync_15_data_out_valid;
  wire                general_fifo_sync_15_data_valid;
  wire                general_fifo_sync_15_full;
  wire                general_fifo_sync_15_empty;
  wire                general_fifo_sync_16_data_in_ready;
  wire       [127:0]  general_fifo_sync_16_data_out;
  wire                general_fifo_sync_16_data_out_valid;
  wire                general_fifo_sync_16_data_valid;
  wire                general_fifo_sync_16_full;
  wire                general_fifo_sync_16_empty;
  wire                general_fifo_sync_17_data_in_ready;
  wire       [127:0]  general_fifo_sync_17_data_out;
  wire                general_fifo_sync_17_data_out_valid;
  wire                general_fifo_sync_17_data_valid;
  wire                general_fifo_sync_17_full;
  wire                general_fifo_sync_17_empty;
  wire                general_fifo_sync_18_data_in_ready;
  wire       [127:0]  general_fifo_sync_18_data_out;
  wire                general_fifo_sync_18_data_out_valid;
  wire                general_fifo_sync_18_data_valid;
  wire                general_fifo_sync_18_full;
  wire                general_fifo_sync_18_empty;
  wire       [1151:0] Configurable_RAM_Norm_doutb;
  wire       [19:0]   mul_add_simd_128_dataOut;
  wire       [19:0]   mul_add_simd_129_dataOut;
  wire       [19:0]   mul_add_simd_130_dataOut;
  wire       [19:0]   mul_add_simd_131_dataOut;
  wire       [19:0]   mul_add_simd_132_dataOut;
  wire       [19:0]   mul_add_simd_133_dataOut;
  wire       [19:0]   mul_add_simd_134_dataOut;
  wire       [19:0]   mul_add_simd_135_dataOut;
  wire       [19:0]   mul_add_simd_136_dataOut;
  wire       [19:0]   mul_add_simd_137_dataOut;
  wire       [19:0]   mul_add_simd_138_dataOut;
  wire       [19:0]   mul_add_simd_139_dataOut;
  wire       [19:0]   mul_add_simd_140_dataOut;
  wire       [19:0]   mul_add_simd_141_dataOut;
  wire       [19:0]   mul_add_simd_142_dataOut;
  wire       [19:0]   mul_add_simd_143_dataOut;
  wire       [19:0]   mul_add_simd_144_dataOut;
  wire       [19:0]   mul_add_simd_145_dataOut;
  wire       [19:0]   mul_add_simd_146_dataOut;
  wire       [19:0]   mul_add_simd_147_dataOut;
  wire       [19:0]   mul_add_simd_148_dataOut;
  wire       [19:0]   mul_add_simd_149_dataOut;
  wire       [19:0]   mul_add_simd_150_dataOut;
  wire       [19:0]   mul_add_simd_151_dataOut;
  wire       [19:0]   mul_add_simd_152_dataOut;
  wire       [19:0]   mul_add_simd_153_dataOut;
  wire       [19:0]   mul_add_simd_154_dataOut;
  wire       [19:0]   mul_add_simd_155_dataOut;
  wire       [19:0]   mul_add_simd_156_dataOut;
  wire       [19:0]   mul_add_simd_157_dataOut;
  wire       [19:0]   mul_add_simd_158_dataOut;
  wire       [19:0]   mul_add_simd_159_dataOut;
  wire       [19:0]   mul_add_simd_160_dataOut;
  wire       [19:0]   mul_add_simd_161_dataOut;
  wire       [19:0]   mul_add_simd_162_dataOut;
  wire       [19:0]   mul_add_simd_163_dataOut;
  wire       [19:0]   mul_add_simd_164_dataOut;
  wire       [19:0]   mul_add_simd_165_dataOut;
  wire       [19:0]   mul_add_simd_166_dataOut;
  wire       [19:0]   mul_add_simd_167_dataOut;
  wire       [19:0]   mul_add_simd_168_dataOut;
  wire       [19:0]   mul_add_simd_169_dataOut;
  wire       [19:0]   mul_add_simd_170_dataOut;
  wire       [19:0]   mul_add_simd_171_dataOut;
  wire       [19:0]   mul_add_simd_172_dataOut;
  wire       [19:0]   mul_add_simd_173_dataOut;
  wire       [19:0]   mul_add_simd_174_dataOut;
  wire       [19:0]   mul_add_simd_175_dataOut;
  wire       [19:0]   mul_add_simd_176_dataOut;
  wire       [19:0]   mul_add_simd_177_dataOut;
  wire       [19:0]   mul_add_simd_178_dataOut;
  wire       [19:0]   mul_add_simd_179_dataOut;
  wire       [19:0]   mul_add_simd_180_dataOut;
  wire       [19:0]   mul_add_simd_181_dataOut;
  wire       [19:0]   mul_add_simd_182_dataOut;
  wire       [19:0]   mul_add_simd_183_dataOut;
  wire       [19:0]   mul_add_simd_184_dataOut;
  wire       [19:0]   mul_add_simd_185_dataOut;
  wire       [19:0]   mul_add_simd_186_dataOut;
  wire       [19:0]   mul_add_simd_187_dataOut;
  wire       [19:0]   mul_add_simd_188_dataOut;
  wire       [19:0]   mul_add_simd_189_dataOut;
  wire       [19:0]   mul_add_simd_190_dataOut;
  wire       [19:0]   mul_add_simd_191_dataOut;
  wire       [19:0]   mul_add_simd_192_dataOut;
  wire       [19:0]   mul_add_simd_193_dataOut;
  wire       [19:0]   mul_add_simd_194_dataOut;
  wire       [19:0]   mul_add_simd_195_dataOut;
  wire       [19:0]   mul_add_simd_196_dataOut;
  wire       [19:0]   mul_add_simd_197_dataOut;
  wire       [19:0]   mul_add_simd_198_dataOut;
  wire       [19:0]   mul_add_simd_199_dataOut;
  wire       [19:0]   mul_add_simd_200_dataOut;
  wire       [19:0]   mul_add_simd_201_dataOut;
  wire       [19:0]   mul_add_simd_202_dataOut;
  wire       [19:0]   mul_add_simd_203_dataOut;
  wire       [19:0]   mul_add_simd_204_dataOut;
  wire       [19:0]   mul_add_simd_205_dataOut;
  wire       [19:0]   mul_add_simd_206_dataOut;
  wire       [19:0]   mul_add_simd_207_dataOut;
  wire       [19:0]   mul_add_simd_208_dataOut;
  wire       [19:0]   mul_add_simd_209_dataOut;
  wire       [19:0]   mul_add_simd_210_dataOut;
  wire       [19:0]   mul_add_simd_211_dataOut;
  wire       [19:0]   mul_add_simd_212_dataOut;
  wire       [19:0]   mul_add_simd_213_dataOut;
  wire       [19:0]   mul_add_simd_214_dataOut;
  wire       [19:0]   mul_add_simd_215_dataOut;
  wire       [19:0]   mul_add_simd_216_dataOut;
  wire       [19:0]   mul_add_simd_217_dataOut;
  wire       [19:0]   mul_add_simd_218_dataOut;
  wire       [19:0]   mul_add_simd_219_dataOut;
  wire       [19:0]   mul_add_simd_220_dataOut;
  wire       [19:0]   mul_add_simd_221_dataOut;
  wire       [19:0]   mul_add_simd_222_dataOut;
  wire       [19:0]   mul_add_simd_223_dataOut;
  wire       [19:0]   mul_add_simd_224_dataOut;
  wire       [19:0]   mul_add_simd_225_dataOut;
  wire       [19:0]   mul_add_simd_226_dataOut;
  wire       [19:0]   mul_add_simd_227_dataOut;
  wire       [19:0]   mul_add_simd_228_dataOut;
  wire       [19:0]   mul_add_simd_229_dataOut;
  wire       [19:0]   mul_add_simd_230_dataOut;
  wire       [19:0]   mul_add_simd_231_dataOut;
  wire       [19:0]   mul_add_simd_232_dataOut;
  wire       [19:0]   mul_add_simd_233_dataOut;
  wire       [19:0]   mul_add_simd_234_dataOut;
  wire       [19:0]   mul_add_simd_235_dataOut;
  wire       [19:0]   mul_add_simd_236_dataOut;
  wire       [19:0]   mul_add_simd_237_dataOut;
  wire       [19:0]   mul_add_simd_238_dataOut;
  wire       [19:0]   mul_add_simd_239_dataOut;
  wire       [19:0]   mul_add_simd_240_dataOut;
  wire       [19:0]   mul_add_simd_241_dataOut;
  wire       [19:0]   mul_add_simd_242_dataOut;
  wire       [19:0]   mul_add_simd_243_dataOut;
  wire       [19:0]   mul_add_simd_244_dataOut;
  wire       [19:0]   mul_add_simd_245_dataOut;
  wire       [19:0]   mul_add_simd_246_dataOut;
  wire       [19:0]   mul_add_simd_247_dataOut;
  wire       [19:0]   mul_add_simd_248_dataOut;
  wire       [19:0]   mul_add_simd_249_dataOut;
  wire       [19:0]   mul_add_simd_250_dataOut;
  wire       [19:0]   mul_add_simd_251_dataOut;
  wire       [19:0]   mul_add_simd_252_dataOut;
  wire       [19:0]   mul_add_simd_253_dataOut;
  wire       [19:0]   mul_add_simd_254_dataOut;
  wire       [19:0]   mul_add_simd_255_dataOut;
  wire       [31:0]   channel_in_acc_8_data_out;
  wire       [31:0]   channel_in_acc_9_data_out;
  wire       [31:0]   channel_in_acc_10_data_out;
  wire       [31:0]   channel_in_acc_11_data_out;
  wire       [31:0]   channel_in_acc_12_data_out;
  wire       [31:0]   channel_in_acc_13_data_out;
  wire       [31:0]   channel_in_acc_14_data_out;
  wire       [31:0]   channel_in_acc_15_data_out;
  wire       [31:0]   channel_out_acc_8_data_out;
  wire       [31:0]   channel_out_acc_9_data_out;
  wire       [31:0]   channel_out_acc_10_data_out;
  wire       [31:0]   channel_out_acc_11_data_out;
  wire       [31:0]   channel_out_acc_12_data_out;
  wire       [31:0]   channel_out_acc_13_data_out;
  wire       [31:0]   channel_out_acc_14_data_out;
  wire       [31:0]   channel_out_acc_15_data_out;
  wire       [5:0]    COMPUTE_TIMES_CHANNEL_IN_REG;
  wire       [7:0]    COMPUTE_TIMES_CHANNEL_IN_REG_8;
  wire       [6:0]    COMPUTE_TIMES_CHANNEL_OUT_REG;
  reg                 compute_ctrl_1_M_Valid_regNext;
  reg        [1151:0] data_fifo_out;
  reg        [127:0]  _zz_data_fifo_out;
  reg        [127:0]  _zz_data_fifo_out_1;
  reg        [127:0]  _zz_data_fifo_out_2;
  reg        [127:0]  _zz_data_fifo_out_3;
  reg        [127:0]  _zz_data_fifo_out_4;
  reg        [127:0]  _zz_data_fifo_out_5;
  reg        [127:0]  _zz_data_fifo_out_6;
  reg        [127:0]  _zz_data_fifo_out_7;
  reg        [127:0]  _zz_data_fifo_out_8;
  wire       [1151:0] ram_temp_output_data;
  reg        [1151:0] ram_temp_output_data_delay_1;
  reg        [1151:0] ram_temp_output_data_delay;
  reg        [71:0]   compute_data_in_0;
  reg        [71:0]   compute_data_in_1;
  reg        [71:0]   compute_data_in_2;
  reg        [71:0]   compute_data_in_3;
  reg        [71:0]   compute_data_in_4;
  reg        [71:0]   compute_data_in_5;
  reg        [71:0]   compute_data_in_6;
  reg        [71:0]   compute_data_in_7;
  reg        [71:0]   compute_data_in_8;
  reg        [71:0]   compute_data_in_9;
  reg        [71:0]   compute_data_in_10;
  reg        [71:0]   compute_data_in_11;
  reg        [71:0]   compute_data_in_12;
  reg        [71:0]   compute_data_in_13;
  reg        [71:0]   compute_data_in_14;
  reg        [71:0]   compute_data_in_15;
  reg        [1151:0] compute_weight_in_0;
  reg        [1151:0] compute_weight_in_1;
  reg        [1151:0] compute_weight_in_2;
  reg        [1151:0] compute_weight_in_3;
  reg        [1151:0] compute_weight_in_4;
  reg        [1151:0] compute_weight_in_5;
  reg        [1151:0] compute_weight_in_6;
  reg        [1151:0] compute_weight_in_7;
  wire       [1151:0] compute_weight_in_delay_0;
  wire       [1151:0] compute_weight_in_delay_1;
  wire       [1151:0] compute_weight_in_delay_2;
  wire       [1151:0] compute_weight_in_delay_3;
  wire       [1151:0] compute_weight_in_delay_4;
  wire       [1151:0] compute_weight_in_delay_5;
  wire       [1151:0] compute_weight_in_delay_6;
  wire       [1151:0] compute_weight_in_delay_7;
  reg        [1151:0] compute_weight_in_0_regNext;
  reg        [1151:0] compute_weight_in_1_regNext;
  reg        [1151:0] compute_weight_in_2_regNext;
  reg        [1151:0] compute_weight_in_3_regNext;
  reg        [1151:0] compute_weight_in_4_regNext;
  reg        [1151:0] compute_weight_in_5_regNext;
  reg        [1151:0] compute_weight_in_6_regNext;
  reg        [1151:0] compute_weight_in_7_regNext;
  reg        [319:0]  compute_data_out_0;
  reg        [319:0]  compute_data_out_1;
  reg        [319:0]  compute_data_out_2;
  reg        [319:0]  compute_data_out_3;
  reg        [319:0]  compute_data_out_4;
  reg        [319:0]  compute_data_out_5;
  reg        [319:0]  compute_data_out_6;
  reg        [319:0]  compute_data_out_7;
  wire       [31:0]   data_result_temp_0;
  wire       [31:0]   data_result_temp_1;
  wire       [31:0]   data_result_temp_2;
  wire       [31:0]   data_result_temp_3;
  wire       [31:0]   data_result_temp_4;
  wire       [31:0]   data_result_temp_5;
  wire       [31:0]   data_result_temp_6;
  wire       [31:0]   data_result_temp_7;

  compute_ctrl compute_ctrl_1 (
    .Start_Cu                          (Start_Cu                                       ), //i
    .Compute_Complete                  (compute_ctrl_1_Compute_Complete                ), //o
    .First_Compute_Complete            (compute_ctrl_1_First_Compute_Complete          ), //o
    .compute_fifo_ready                (compute_ctrl_1_compute_fifo_ready              ), //i
    .rd_en_fifo                        (compute_ctrl_1_rd_en_fifo                      ), //o
    .M_ready                           (M_DATA_ready                                   ), //i
    .M_Valid                           (compute_ctrl_1_M_Valid                         ), //o
    .weight_addrb                      (compute_ctrl_1_weight_addrb                    ), //o
    .ram_temp_read_address             (compute_ctrl_1_ram_temp_read_address           ), //o
    .ram_temp_write_address            (compute_ctrl_1_ram_temp_write_address          ), //o
    .COMPUTE_TIMES_CHANNEL_IN_REG      (compute_ctrl_1_COMPUTE_TIMES_CHANNEL_IN_REG    ), //i
    .COMPUTE_TIMES_CHANNEL_IN_REG_8    (compute_ctrl_1_COMPUTE_TIMES_CHANNEL_IN_REG_8  ), //i
    .COMPUTE_TIMES_CHANNEL_OUT_REG     (compute_ctrl_1_COMPUTE_TIMES_CHANNEL_OUT_REG   ), //i
    .ROW_NUM_CHANNEL_OUT_REG           (Row_Num_Out_REG                                ), //i
    .S_Count_Fifo                      (compute_ctrl_1_S_Count_Fifo                    ), //o
    .M_Count_Fifo                      (compute_ctrl_1_M_Count_Fifo                    ), //o
    .clk                               (clk                                            ), //i
    .reset                             (reset                                          )  //i
  );
  load_weight load_weight_1 (
    .Start_Pa                 (Start_Pa                            ), //i
    .Weight_Single_Num_REG    (Weight_Single_Num_REG               ), //i
    .Bias_Num_REG             (Bias_Num_REG                        ), //i
    .Write_Block_Complete     (load_weight_1_Write_Block_Complete  ), //o
    .S_Para_Data_valid        (para_data_valid                     ), //i
    .S_Para_Data_ready        (load_weight_1_S_Para_Data_ready     ), //o
    .S_Para_Data_payload      (para_data_payload                   ), //i
    .Weight_Addrb             (compute_ctrl_1_weight_addrb         ), //i
    .Data_Out_Weight_0        (load_weight_1_Data_Out_Weight_0     ), //o
    .Data_Out_Weight_1        (load_weight_1_Data_Out_Weight_1     ), //o
    .Data_Out_Weight_2        (load_weight_1_Data_Out_Weight_2     ), //o
    .Data_Out_Weight_3        (load_weight_1_Data_Out_Weight_3     ), //o
    .Data_Out_Weight_4        (load_weight_1_Data_Out_Weight_4     ), //o
    .Data_Out_Weight_5        (load_weight_1_Data_Out_Weight_5     ), //o
    .Data_Out_Weight_6        (load_weight_1_Data_Out_Weight_6     ), //o
    .Data_Out_Weight_7        (load_weight_1_Data_Out_Weight_7     ), //o
    .Data_Out_Weight_8        (load_weight_1_Data_Out_Weight_8     ), //o
    .Bias_Addrb               (Bias_Addrb                          ), //i
    .Data_Out_Bias            (load_weight_1_Data_Out_Bias         ), //o
    .Data_Out_Scale           (load_weight_1_Data_Out_Scale        ), //o
    .Data_Out_Shift           (load_weight_1_Data_Out_Shift        ), //o
    .clk                      (clk                                 ), //i
    .reset                    (reset                               )  //i
  );
  general_fifo_sync_1 general_fifo_sync_10 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_10_data_in         ), //i
    .wr_en             (general_fifo_sync_10_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_10_data_in_ready   ), //o
    .data_out          (general_fifo_sync_10_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_10_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_10_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_10_s_data_count    ), //i
    .data_valid        (general_fifo_sync_10_data_valid      ), //o
    .full              (general_fifo_sync_10_full            ), //o
    .empty             (general_fifo_sync_10_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_11 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_11_data_in         ), //i
    .wr_en             (general_fifo_sync_11_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_11_data_in_ready   ), //o
    .data_out          (general_fifo_sync_11_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_11_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_11_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_11_s_data_count    ), //i
    .data_valid        (general_fifo_sync_11_data_valid      ), //o
    .full              (general_fifo_sync_11_full            ), //o
    .empty             (general_fifo_sync_11_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_12 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_12_data_in         ), //i
    .wr_en             (general_fifo_sync_12_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_12_data_in_ready   ), //o
    .data_out          (general_fifo_sync_12_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_12_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_12_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_12_s_data_count    ), //i
    .data_valid        (general_fifo_sync_12_data_valid      ), //o
    .full              (general_fifo_sync_12_full            ), //o
    .empty             (general_fifo_sync_12_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_13 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_13_data_in         ), //i
    .wr_en             (general_fifo_sync_13_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_13_data_in_ready   ), //o
    .data_out          (general_fifo_sync_13_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_13_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_13_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_13_s_data_count    ), //i
    .data_valid        (general_fifo_sync_13_data_valid      ), //o
    .full              (general_fifo_sync_13_full            ), //o
    .empty             (general_fifo_sync_13_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_14 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_14_data_in         ), //i
    .wr_en             (general_fifo_sync_14_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_14_data_in_ready   ), //o
    .data_out          (general_fifo_sync_14_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_14_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_14_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_14_s_data_count    ), //i
    .data_valid        (general_fifo_sync_14_data_valid      ), //o
    .full              (general_fifo_sync_14_full            ), //o
    .empty             (general_fifo_sync_14_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_15 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_15_data_in         ), //i
    .wr_en             (general_fifo_sync_15_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_15_data_in_ready   ), //o
    .data_out          (general_fifo_sync_15_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_15_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_15_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_15_s_data_count    ), //i
    .data_valid        (general_fifo_sync_15_data_valid      ), //o
    .full              (general_fifo_sync_15_full            ), //o
    .empty             (general_fifo_sync_15_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_16 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_16_data_in         ), //i
    .wr_en             (general_fifo_sync_16_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_16_data_in_ready   ), //o
    .data_out          (general_fifo_sync_16_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_16_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_16_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_16_s_data_count    ), //i
    .data_valid        (general_fifo_sync_16_data_valid      ), //o
    .full              (general_fifo_sync_16_full            ), //o
    .empty             (general_fifo_sync_16_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_17 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_17_data_in         ), //i
    .wr_en             (general_fifo_sync_17_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_17_data_in_ready   ), //o
    .data_out          (general_fifo_sync_17_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_17_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_17_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_17_s_data_count    ), //i
    .data_valid        (general_fifo_sync_17_data_valid      ), //o
    .full              (general_fifo_sync_17_full            ), //o
    .empty             (general_fifo_sync_17_empty           )  //o
  );
  general_fifo_sync_1 general_fifo_sync_18 (
    .reset             (reset                                ), //i
    .clk               (clk                                  ), //i
    .data_in           (general_fifo_sync_18_data_in         ), //i
    .wr_en             (general_fifo_sync_18_wr_en           ), //i
    .data_in_ready     (general_fifo_sync_18_data_in_ready   ), //o
    .data_out          (general_fifo_sync_18_data_out        ), //o
    .rd_en             (compute_ctrl_1_rd_en_fifo            ), //i
    .data_out_valid    (general_fifo_sync_18_data_out_valid  ), //o
    .m_data_count      (general_fifo_sync_18_m_data_count    ), //i
    .s_data_count      (general_fifo_sync_18_s_data_count    ), //i
    .data_valid        (general_fifo_sync_18_data_valid      ), //o
    .full              (general_fifo_sync_18_full            ), //o
    .empty             (general_fifo_sync_18_empty           )  //o
  );
  sdpram_16 Configurable_RAM_Norm (
    .doutb    (Configurable_RAM_Norm_doutb            ), //o
    .addra    (compute_ctrl_1_ram_temp_write_address  ), //i
    .addrb    (compute_ctrl_1_ram_temp_read_address   ), //i
    .dina     (data_fifo_out                          ), //i
    .ena      (1'b1                                   ), //i
    .enb      (1'b1                                   ), //i
    .wea      (Configurable_RAM_Norm_wea              ), //i
    .clk      (clk                                    )  //i
  );
  mul_add_simd mul_add_simd_128 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_128_weightIn  ), //i
    .dataOut     (mul_add_simd_128_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_129 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_129_weightIn  ), //i
    .dataOut     (mul_add_simd_129_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_130 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_130_weightIn  ), //i
    .dataOut     (mul_add_simd_130_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_131 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_131_weightIn  ), //i
    .dataOut     (mul_add_simd_131_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_132 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_132_weightIn  ), //i
    .dataOut     (mul_add_simd_132_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_133 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_133_weightIn  ), //i
    .dataOut     (mul_add_simd_133_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_134 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_134_weightIn  ), //i
    .dataOut     (mul_add_simd_134_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_135 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_135_weightIn  ), //i
    .dataOut     (mul_add_simd_135_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_136 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_136_weightIn  ), //i
    .dataOut     (mul_add_simd_136_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_137 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_137_weightIn  ), //i
    .dataOut     (mul_add_simd_137_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_138 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_138_weightIn  ), //i
    .dataOut     (mul_add_simd_138_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_139 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_139_weightIn  ), //i
    .dataOut     (mul_add_simd_139_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_140 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_140_weightIn  ), //i
    .dataOut     (mul_add_simd_140_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_141 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_141_weightIn  ), //i
    .dataOut     (mul_add_simd_141_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_142 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_142_weightIn  ), //i
    .dataOut     (mul_add_simd_142_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_143 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_143_weightIn  ), //i
    .dataOut     (mul_add_simd_143_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_144 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_144_weightIn  ), //i
    .dataOut     (mul_add_simd_144_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_145 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_145_weightIn  ), //i
    .dataOut     (mul_add_simd_145_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_146 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_146_weightIn  ), //i
    .dataOut     (mul_add_simd_146_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_147 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_147_weightIn  ), //i
    .dataOut     (mul_add_simd_147_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_148 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_148_weightIn  ), //i
    .dataOut     (mul_add_simd_148_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_149 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_149_weightIn  ), //i
    .dataOut     (mul_add_simd_149_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_150 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_150_weightIn  ), //i
    .dataOut     (mul_add_simd_150_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_151 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_151_weightIn  ), //i
    .dataOut     (mul_add_simd_151_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_152 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_152_weightIn  ), //i
    .dataOut     (mul_add_simd_152_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_153 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_153_weightIn  ), //i
    .dataOut     (mul_add_simd_153_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_154 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_154_weightIn  ), //i
    .dataOut     (mul_add_simd_154_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_155 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_155_weightIn  ), //i
    .dataOut     (mul_add_simd_155_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_156 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_156_weightIn  ), //i
    .dataOut     (mul_add_simd_156_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_157 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_157_weightIn  ), //i
    .dataOut     (mul_add_simd_157_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_158 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_158_weightIn  ), //i
    .dataOut     (mul_add_simd_158_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_159 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_159_weightIn  ), //i
    .dataOut     (mul_add_simd_159_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_160 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_160_weightIn  ), //i
    .dataOut     (mul_add_simd_160_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_161 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_161_weightIn  ), //i
    .dataOut     (mul_add_simd_161_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_162 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_162_weightIn  ), //i
    .dataOut     (mul_add_simd_162_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_163 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_163_weightIn  ), //i
    .dataOut     (mul_add_simd_163_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_164 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_164_weightIn  ), //i
    .dataOut     (mul_add_simd_164_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_165 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_165_weightIn  ), //i
    .dataOut     (mul_add_simd_165_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_166 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_166_weightIn  ), //i
    .dataOut     (mul_add_simd_166_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_167 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_167_weightIn  ), //i
    .dataOut     (mul_add_simd_167_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_168 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_168_weightIn  ), //i
    .dataOut     (mul_add_simd_168_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_169 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_169_weightIn  ), //i
    .dataOut     (mul_add_simd_169_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_170 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_170_weightIn  ), //i
    .dataOut     (mul_add_simd_170_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_171 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_171_weightIn  ), //i
    .dataOut     (mul_add_simd_171_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_172 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_172_weightIn  ), //i
    .dataOut     (mul_add_simd_172_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_173 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_173_weightIn  ), //i
    .dataOut     (mul_add_simd_173_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_174 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_174_weightIn  ), //i
    .dataOut     (mul_add_simd_174_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_175 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_175_weightIn  ), //i
    .dataOut     (mul_add_simd_175_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_176 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_176_weightIn  ), //i
    .dataOut     (mul_add_simd_176_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_177 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_177_weightIn  ), //i
    .dataOut     (mul_add_simd_177_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_178 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_178_weightIn  ), //i
    .dataOut     (mul_add_simd_178_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_179 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_179_weightIn  ), //i
    .dataOut     (mul_add_simd_179_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_180 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_180_weightIn  ), //i
    .dataOut     (mul_add_simd_180_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_181 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_181_weightIn  ), //i
    .dataOut     (mul_add_simd_181_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_182 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_182_weightIn  ), //i
    .dataOut     (mul_add_simd_182_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_183 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_183_weightIn  ), //i
    .dataOut     (mul_add_simd_183_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_184 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_184_weightIn  ), //i
    .dataOut     (mul_add_simd_184_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_185 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_185_weightIn  ), //i
    .dataOut     (mul_add_simd_185_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_186 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_186_weightIn  ), //i
    .dataOut     (mul_add_simd_186_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_187 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_187_weightIn  ), //i
    .dataOut     (mul_add_simd_187_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_188 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_188_weightIn  ), //i
    .dataOut     (mul_add_simd_188_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_189 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_189_weightIn  ), //i
    .dataOut     (mul_add_simd_189_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_190 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_190_weightIn  ), //i
    .dataOut     (mul_add_simd_190_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_191 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_191_weightIn  ), //i
    .dataOut     (mul_add_simd_191_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_192 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_192_weightIn  ), //i
    .dataOut     (mul_add_simd_192_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_193 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_193_weightIn  ), //i
    .dataOut     (mul_add_simd_193_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_194 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_194_weightIn  ), //i
    .dataOut     (mul_add_simd_194_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_195 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_195_weightIn  ), //i
    .dataOut     (mul_add_simd_195_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_196 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_196_weightIn  ), //i
    .dataOut     (mul_add_simd_196_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_197 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_197_weightIn  ), //i
    .dataOut     (mul_add_simd_197_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_198 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_198_weightIn  ), //i
    .dataOut     (mul_add_simd_198_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_199 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_199_weightIn  ), //i
    .dataOut     (mul_add_simd_199_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_200 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_200_weightIn  ), //i
    .dataOut     (mul_add_simd_200_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_201 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_201_weightIn  ), //i
    .dataOut     (mul_add_simd_201_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_202 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_202_weightIn  ), //i
    .dataOut     (mul_add_simd_202_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_203 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_203_weightIn  ), //i
    .dataOut     (mul_add_simd_203_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_204 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_204_weightIn  ), //i
    .dataOut     (mul_add_simd_204_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_205 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_205_weightIn  ), //i
    .dataOut     (mul_add_simd_205_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_206 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_206_weightIn  ), //i
    .dataOut     (mul_add_simd_206_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_207 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_207_weightIn  ), //i
    .dataOut     (mul_add_simd_207_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_208 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_208_weightIn  ), //i
    .dataOut     (mul_add_simd_208_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_209 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_209_weightIn  ), //i
    .dataOut     (mul_add_simd_209_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_210 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_210_weightIn  ), //i
    .dataOut     (mul_add_simd_210_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_211 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_211_weightIn  ), //i
    .dataOut     (mul_add_simd_211_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_212 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_212_weightIn  ), //i
    .dataOut     (mul_add_simd_212_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_213 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_213_weightIn  ), //i
    .dataOut     (mul_add_simd_213_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_214 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_214_weightIn  ), //i
    .dataOut     (mul_add_simd_214_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_215 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_215_weightIn  ), //i
    .dataOut     (mul_add_simd_215_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_216 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_216_weightIn  ), //i
    .dataOut     (mul_add_simd_216_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_217 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_217_weightIn  ), //i
    .dataOut     (mul_add_simd_217_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_218 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_218_weightIn  ), //i
    .dataOut     (mul_add_simd_218_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_219 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_219_weightIn  ), //i
    .dataOut     (mul_add_simd_219_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_220 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_220_weightIn  ), //i
    .dataOut     (mul_add_simd_220_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_221 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_221_weightIn  ), //i
    .dataOut     (mul_add_simd_221_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_222 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_222_weightIn  ), //i
    .dataOut     (mul_add_simd_222_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_223 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_223_weightIn  ), //i
    .dataOut     (mul_add_simd_223_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_224 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_224_weightIn  ), //i
    .dataOut     (mul_add_simd_224_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_225 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_225_weightIn  ), //i
    .dataOut     (mul_add_simd_225_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_226 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_226_weightIn  ), //i
    .dataOut     (mul_add_simd_226_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_227 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_227_weightIn  ), //i
    .dataOut     (mul_add_simd_227_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_228 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_228_weightIn  ), //i
    .dataOut     (mul_add_simd_228_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_229 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_229_weightIn  ), //i
    .dataOut     (mul_add_simd_229_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_230 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_230_weightIn  ), //i
    .dataOut     (mul_add_simd_230_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_231 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_231_weightIn  ), //i
    .dataOut     (mul_add_simd_231_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_232 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_232_weightIn  ), //i
    .dataOut     (mul_add_simd_232_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_233 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_233_weightIn  ), //i
    .dataOut     (mul_add_simd_233_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_234 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_234_weightIn  ), //i
    .dataOut     (mul_add_simd_234_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_235 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_235_weightIn  ), //i
    .dataOut     (mul_add_simd_235_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_236 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_236_weightIn  ), //i
    .dataOut     (mul_add_simd_236_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_237 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_237_weightIn  ), //i
    .dataOut     (mul_add_simd_237_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_238 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_238_weightIn  ), //i
    .dataOut     (mul_add_simd_238_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_239 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_239_weightIn  ), //i
    .dataOut     (mul_add_simd_239_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_240 (
    .dataIn      (compute_data_in_0          ), //i
    .weightIn    (mul_add_simd_240_weightIn  ), //i
    .dataOut     (mul_add_simd_240_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_241 (
    .dataIn      (compute_data_in_1          ), //i
    .weightIn    (mul_add_simd_241_weightIn  ), //i
    .dataOut     (mul_add_simd_241_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_242 (
    .dataIn      (compute_data_in_2          ), //i
    .weightIn    (mul_add_simd_242_weightIn  ), //i
    .dataOut     (mul_add_simd_242_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_243 (
    .dataIn      (compute_data_in_3          ), //i
    .weightIn    (mul_add_simd_243_weightIn  ), //i
    .dataOut     (mul_add_simd_243_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_244 (
    .dataIn      (compute_data_in_4          ), //i
    .weightIn    (mul_add_simd_244_weightIn  ), //i
    .dataOut     (mul_add_simd_244_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_245 (
    .dataIn      (compute_data_in_5          ), //i
    .weightIn    (mul_add_simd_245_weightIn  ), //i
    .dataOut     (mul_add_simd_245_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_246 (
    .dataIn      (compute_data_in_6          ), //i
    .weightIn    (mul_add_simd_246_weightIn  ), //i
    .dataOut     (mul_add_simd_246_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_247 (
    .dataIn      (compute_data_in_7          ), //i
    .weightIn    (mul_add_simd_247_weightIn  ), //i
    .dataOut     (mul_add_simd_247_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_248 (
    .dataIn      (compute_data_in_8          ), //i
    .weightIn    (mul_add_simd_248_weightIn  ), //i
    .dataOut     (mul_add_simd_248_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_249 (
    .dataIn      (compute_data_in_9          ), //i
    .weightIn    (mul_add_simd_249_weightIn  ), //i
    .dataOut     (mul_add_simd_249_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_250 (
    .dataIn      (compute_data_in_10         ), //i
    .weightIn    (mul_add_simd_250_weightIn  ), //i
    .dataOut     (mul_add_simd_250_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_251 (
    .dataIn      (compute_data_in_11         ), //i
    .weightIn    (mul_add_simd_251_weightIn  ), //i
    .dataOut     (mul_add_simd_251_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_252 (
    .dataIn      (compute_data_in_12         ), //i
    .weightIn    (mul_add_simd_252_weightIn  ), //i
    .dataOut     (mul_add_simd_252_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_253 (
    .dataIn      (compute_data_in_13         ), //i
    .weightIn    (mul_add_simd_253_weightIn  ), //i
    .dataOut     (mul_add_simd_253_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_254 (
    .dataIn      (compute_data_in_14         ), //i
    .weightIn    (mul_add_simd_254_weightIn  ), //i
    .dataOut     (mul_add_simd_254_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  mul_add_simd mul_add_simd_255 (
    .dataIn      (compute_data_in_15         ), //i
    .weightIn    (mul_add_simd_255_weightIn  ), //i
    .dataOut     (mul_add_simd_255_dataOut   ), //o
    .clk         (clk                        ), //i
    .reset       (reset                      )  //i
  );
  channel_in_acc channel_in_acc_8 (
    .data_in     (compute_data_out_0         ), //i
    .data_out    (channel_in_acc_8_data_out  ), //o
    .clk         (clk                        )  //i
  );
  channel_in_acc channel_in_acc_9 (
    .data_in     (compute_data_out_1         ), //i
    .data_out    (channel_in_acc_9_data_out  ), //o
    .clk         (clk                        )  //i
  );
  channel_in_acc channel_in_acc_10 (
    .data_in     (compute_data_out_2          ), //i
    .data_out    (channel_in_acc_10_data_out  ), //o
    .clk         (clk                         )  //i
  );
  channel_in_acc channel_in_acc_11 (
    .data_in     (compute_data_out_3          ), //i
    .data_out    (channel_in_acc_11_data_out  ), //o
    .clk         (clk                         )  //i
  );
  channel_in_acc channel_in_acc_12 (
    .data_in     (compute_data_out_4          ), //i
    .data_out    (channel_in_acc_12_data_out  ), //o
    .clk         (clk                         )  //i
  );
  channel_in_acc channel_in_acc_13 (
    .data_in     (compute_data_out_5          ), //i
    .data_out    (channel_in_acc_13_data_out  ), //o
    .clk         (clk                         )  //i
  );
  channel_in_acc channel_in_acc_14 (
    .data_in     (compute_data_out_6          ), //i
    .data_out    (channel_in_acc_14_data_out  ), //o
    .clk         (clk                         )  //i
  );
  channel_in_acc channel_in_acc_15 (
    .data_in     (compute_data_out_7          ), //i
    .data_out    (channel_in_acc_15_data_out  ), //o
    .clk         (clk                         )  //i
  );
  channel_out_acc channel_out_acc_8 (
    .data_in                   (channel_in_acc_8_data_out              ), //i
    .data_out                  (channel_out_acc_8_data_out             ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_9 (
    .data_in                   (channel_in_acc_9_data_out              ), //i
    .data_out                  (channel_out_acc_9_data_out             ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_10 (
    .data_in                   (channel_in_acc_10_data_out             ), //i
    .data_out                  (channel_out_acc_10_data_out            ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_11 (
    .data_in                   (channel_in_acc_11_data_out             ), //i
    .data_out                  (channel_out_acc_11_data_out            ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_12 (
    .data_in                   (channel_in_acc_12_data_out             ), //i
    .data_out                  (channel_out_acc_12_data_out            ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_13 (
    .data_in                   (channel_in_acc_13_data_out             ), //i
    .data_out                  (channel_out_acc_13_data_out            ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_14 (
    .data_in                   (channel_in_acc_14_data_out             ), //i
    .data_out                  (channel_out_acc_14_data_out            ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  channel_out_acc channel_out_acc_15 (
    .data_in                   (channel_in_acc_15_data_out             ), //i
    .data_out                  (channel_out_acc_15_data_out            ), //o
    .First_Compute_Complete    (compute_ctrl_1_First_Compute_Complete  ), //i
    .clk                       (clk                                    ), //i
    .reset                     (reset                                  )  //i
  );
  assign COMPUTE_TIMES_CHANNEL_IN_REG = (Channel_In_Num_REG >>> 4);
  assign COMPUTE_TIMES_CHANNEL_IN_REG_8 = (Channel_In_Num_REG >>> 2);
  assign COMPUTE_TIMES_CHANNEL_OUT_REG = (Channel_Out_Num_REG >>> 3);
  assign compute_ctrl_1_COMPUTE_TIMES_CHANNEL_IN_REG = {5'd0, COMPUTE_TIMES_CHANNEL_IN_REG};
  assign compute_ctrl_1_COMPUTE_TIMES_CHANNEL_IN_REG_8 = {3'd0, COMPUTE_TIMES_CHANNEL_IN_REG_8};
  assign compute_ctrl_1_COMPUTE_TIMES_CHANNEL_OUT_REG = {4'd0, COMPUTE_TIMES_CHANNEL_OUT_REG};
  assign Compute_Complete = compute_ctrl_1_Compute_Complete;
  assign Write_Block_Complete = load_weight_1_Write_Block_Complete;
  assign para_data_ready = load_weight_1_S_Para_Data_ready;
  assign Data_Out_Bias = load_weight_1_Data_Out_Bias;
  assign Data_Out_Scale = load_weight_1_Data_Out_Scale;
  assign Data_Out_Shift = load_weight_1_Data_Out_Shift;
  assign general_fifo_sync_10_wr_en = S_DATA_Valid[0];
  assign general_fifo_sync_10_data_in = S_DATA[63 : 0];
  assign general_fifo_sync_10_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_10_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out[63 : 0] = general_fifo_sync_10_data_out[127 : 64];
    _zz_data_fifo_out[127 : 64] = general_fifo_sync_10_data_out[63 : 0];
  end

  always @(*) begin
    data_fifo_out[127 : 0] = _zz_data_fifo_out;
    data_fifo_out[255 : 128] = _zz_data_fifo_out_1;
    data_fifo_out[383 : 256] = _zz_data_fifo_out_2;
    data_fifo_out[511 : 384] = _zz_data_fifo_out_3;
    data_fifo_out[639 : 512] = _zz_data_fifo_out_4;
    data_fifo_out[767 : 640] = _zz_data_fifo_out_5;
    data_fifo_out[895 : 768] = _zz_data_fifo_out_6;
    data_fifo_out[1023 : 896] = _zz_data_fifo_out_7;
    data_fifo_out[1151 : 1024] = _zz_data_fifo_out_8;
  end

  assign general_fifo_sync_11_wr_en = S_DATA_Valid[1];
  assign general_fifo_sync_11_data_in = S_DATA[127 : 64];
  assign general_fifo_sync_11_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_11_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_1[63 : 0] = general_fifo_sync_11_data_out[127 : 64];
    _zz_data_fifo_out_1[127 : 64] = general_fifo_sync_11_data_out[63 : 0];
  end

  assign general_fifo_sync_12_wr_en = S_DATA_Valid[2];
  assign general_fifo_sync_12_data_in = S_DATA[191 : 128];
  assign general_fifo_sync_12_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_12_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_2[63 : 0] = general_fifo_sync_12_data_out[127 : 64];
    _zz_data_fifo_out_2[127 : 64] = general_fifo_sync_12_data_out[63 : 0];
  end

  assign general_fifo_sync_13_wr_en = S_DATA_Valid[3];
  assign general_fifo_sync_13_data_in = S_DATA[255 : 192];
  assign general_fifo_sync_13_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_13_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_3[63 : 0] = general_fifo_sync_13_data_out[127 : 64];
    _zz_data_fifo_out_3[127 : 64] = general_fifo_sync_13_data_out[63 : 0];
  end

  assign general_fifo_sync_14_wr_en = S_DATA_Valid[4];
  assign general_fifo_sync_14_data_in = S_DATA[319 : 256];
  assign general_fifo_sync_14_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_14_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_4[63 : 0] = general_fifo_sync_14_data_out[127 : 64];
    _zz_data_fifo_out_4[127 : 64] = general_fifo_sync_14_data_out[63 : 0];
  end

  assign general_fifo_sync_15_wr_en = S_DATA_Valid[5];
  assign general_fifo_sync_15_data_in = S_DATA[383 : 320];
  assign general_fifo_sync_15_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_15_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_5[63 : 0] = general_fifo_sync_15_data_out[127 : 64];
    _zz_data_fifo_out_5[127 : 64] = general_fifo_sync_15_data_out[63 : 0];
  end

  assign general_fifo_sync_16_wr_en = S_DATA_Valid[6];
  assign general_fifo_sync_16_data_in = S_DATA[447 : 384];
  assign general_fifo_sync_16_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_16_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_6[63 : 0] = general_fifo_sync_16_data_out[127 : 64];
    _zz_data_fifo_out_6[127 : 64] = general_fifo_sync_16_data_out[63 : 0];
  end

  assign general_fifo_sync_17_wr_en = S_DATA_Valid[7];
  assign general_fifo_sync_17_data_in = S_DATA[511 : 448];
  assign general_fifo_sync_17_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_17_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_7[63 : 0] = general_fifo_sync_17_data_out[127 : 64];
    _zz_data_fifo_out_7[127 : 64] = general_fifo_sync_17_data_out[63 : 0];
  end

  assign general_fifo_sync_18_wr_en = S_DATA_Valid[8];
  assign general_fifo_sync_18_data_in = S_DATA[575 : 512];
  assign general_fifo_sync_18_m_data_count = compute_ctrl_1_M_Count_Fifo;
  assign general_fifo_sync_18_s_data_count = compute_ctrl_1_S_Count_Fifo;
  always @(*) begin
    _zz_data_fifo_out_8[63 : 0] = general_fifo_sync_18_data_out[127 : 64];
    _zz_data_fifo_out_8[127 : 64] = general_fifo_sync_18_data_out[63 : 0];
  end

  assign S_DATA_Ready = ((general_fifo_sync_10_data_in_ready && general_fifo_sync_11_data_in_ready) && general_fifo_sync_12_data_in_ready);
  assign compute_ctrl_1_compute_fifo_ready = ((general_fifo_sync_10_data_out_valid && general_fifo_sync_11_data_out_valid) && general_fifo_sync_12_data_out_valid);
  assign Configurable_RAM_Norm_wea = compute_ctrl_1_rd_en_fifo;
  assign ram_temp_output_data = Configurable_RAM_Norm_doutb;
  always @(*) begin
    compute_data_in_0[7 : 0] = ram_temp_output_data[7 : 0];
    compute_data_in_0[15 : 8] = ram_temp_output_data[135 : 128];
    compute_data_in_0[23 : 16] = ram_temp_output_data[263 : 256];
    compute_data_in_0[31 : 24] = ram_temp_output_data[391 : 384];
    compute_data_in_0[39 : 32] = ram_temp_output_data[519 : 512];
    compute_data_in_0[47 : 40] = ram_temp_output_data[647 : 640];
    compute_data_in_0[55 : 48] = ram_temp_output_data[775 : 768];
    compute_data_in_0[63 : 56] = ram_temp_output_data[903 : 896];
    compute_data_in_0[71 : 64] = ram_temp_output_data[1031 : 1024];
  end

  always @(*) begin
    compute_data_in_1[7 : 0] = ram_temp_output_data[15 : 8];
    compute_data_in_1[15 : 8] = ram_temp_output_data[143 : 136];
    compute_data_in_1[23 : 16] = ram_temp_output_data[271 : 264];
    compute_data_in_1[31 : 24] = ram_temp_output_data[399 : 392];
    compute_data_in_1[39 : 32] = ram_temp_output_data[527 : 520];
    compute_data_in_1[47 : 40] = ram_temp_output_data[655 : 648];
    compute_data_in_1[55 : 48] = ram_temp_output_data[783 : 776];
    compute_data_in_1[63 : 56] = ram_temp_output_data[911 : 904];
    compute_data_in_1[71 : 64] = ram_temp_output_data[1039 : 1032];
  end

  always @(*) begin
    compute_data_in_2[7 : 0] = ram_temp_output_data[23 : 16];
    compute_data_in_2[15 : 8] = ram_temp_output_data[151 : 144];
    compute_data_in_2[23 : 16] = ram_temp_output_data[279 : 272];
    compute_data_in_2[31 : 24] = ram_temp_output_data[407 : 400];
    compute_data_in_2[39 : 32] = ram_temp_output_data[535 : 528];
    compute_data_in_2[47 : 40] = ram_temp_output_data[663 : 656];
    compute_data_in_2[55 : 48] = ram_temp_output_data[791 : 784];
    compute_data_in_2[63 : 56] = ram_temp_output_data[919 : 912];
    compute_data_in_2[71 : 64] = ram_temp_output_data[1047 : 1040];
  end

  always @(*) begin
    compute_data_in_3[7 : 0] = ram_temp_output_data[31 : 24];
    compute_data_in_3[15 : 8] = ram_temp_output_data[159 : 152];
    compute_data_in_3[23 : 16] = ram_temp_output_data[287 : 280];
    compute_data_in_3[31 : 24] = ram_temp_output_data[415 : 408];
    compute_data_in_3[39 : 32] = ram_temp_output_data[543 : 536];
    compute_data_in_3[47 : 40] = ram_temp_output_data[671 : 664];
    compute_data_in_3[55 : 48] = ram_temp_output_data[799 : 792];
    compute_data_in_3[63 : 56] = ram_temp_output_data[927 : 920];
    compute_data_in_3[71 : 64] = ram_temp_output_data[1055 : 1048];
  end

  always @(*) begin
    compute_data_in_4[7 : 0] = ram_temp_output_data[39 : 32];
    compute_data_in_4[15 : 8] = ram_temp_output_data[167 : 160];
    compute_data_in_4[23 : 16] = ram_temp_output_data[295 : 288];
    compute_data_in_4[31 : 24] = ram_temp_output_data[423 : 416];
    compute_data_in_4[39 : 32] = ram_temp_output_data[551 : 544];
    compute_data_in_4[47 : 40] = ram_temp_output_data[679 : 672];
    compute_data_in_4[55 : 48] = ram_temp_output_data[807 : 800];
    compute_data_in_4[63 : 56] = ram_temp_output_data[935 : 928];
    compute_data_in_4[71 : 64] = ram_temp_output_data[1063 : 1056];
  end

  always @(*) begin
    compute_data_in_5[7 : 0] = ram_temp_output_data[47 : 40];
    compute_data_in_5[15 : 8] = ram_temp_output_data[175 : 168];
    compute_data_in_5[23 : 16] = ram_temp_output_data[303 : 296];
    compute_data_in_5[31 : 24] = ram_temp_output_data[431 : 424];
    compute_data_in_5[39 : 32] = ram_temp_output_data[559 : 552];
    compute_data_in_5[47 : 40] = ram_temp_output_data[687 : 680];
    compute_data_in_5[55 : 48] = ram_temp_output_data[815 : 808];
    compute_data_in_5[63 : 56] = ram_temp_output_data[943 : 936];
    compute_data_in_5[71 : 64] = ram_temp_output_data[1071 : 1064];
  end

  always @(*) begin
    compute_data_in_6[7 : 0] = ram_temp_output_data[55 : 48];
    compute_data_in_6[15 : 8] = ram_temp_output_data[183 : 176];
    compute_data_in_6[23 : 16] = ram_temp_output_data[311 : 304];
    compute_data_in_6[31 : 24] = ram_temp_output_data[439 : 432];
    compute_data_in_6[39 : 32] = ram_temp_output_data[567 : 560];
    compute_data_in_6[47 : 40] = ram_temp_output_data[695 : 688];
    compute_data_in_6[55 : 48] = ram_temp_output_data[823 : 816];
    compute_data_in_6[63 : 56] = ram_temp_output_data[951 : 944];
    compute_data_in_6[71 : 64] = ram_temp_output_data[1079 : 1072];
  end

  always @(*) begin
    compute_data_in_7[7 : 0] = ram_temp_output_data[63 : 56];
    compute_data_in_7[15 : 8] = ram_temp_output_data[191 : 184];
    compute_data_in_7[23 : 16] = ram_temp_output_data[319 : 312];
    compute_data_in_7[31 : 24] = ram_temp_output_data[447 : 440];
    compute_data_in_7[39 : 32] = ram_temp_output_data[575 : 568];
    compute_data_in_7[47 : 40] = ram_temp_output_data[703 : 696];
    compute_data_in_7[55 : 48] = ram_temp_output_data[831 : 824];
    compute_data_in_7[63 : 56] = ram_temp_output_data[959 : 952];
    compute_data_in_7[71 : 64] = ram_temp_output_data[1087 : 1080];
  end

  always @(*) begin
    compute_data_in_8[7 : 0] = ram_temp_output_data[71 : 64];
    compute_data_in_8[15 : 8] = ram_temp_output_data[199 : 192];
    compute_data_in_8[23 : 16] = ram_temp_output_data[327 : 320];
    compute_data_in_8[31 : 24] = ram_temp_output_data[455 : 448];
    compute_data_in_8[39 : 32] = ram_temp_output_data[583 : 576];
    compute_data_in_8[47 : 40] = ram_temp_output_data[711 : 704];
    compute_data_in_8[55 : 48] = ram_temp_output_data[839 : 832];
    compute_data_in_8[63 : 56] = ram_temp_output_data[967 : 960];
    compute_data_in_8[71 : 64] = ram_temp_output_data[1095 : 1088];
  end

  always @(*) begin
    compute_data_in_9[7 : 0] = ram_temp_output_data[79 : 72];
    compute_data_in_9[15 : 8] = ram_temp_output_data[207 : 200];
    compute_data_in_9[23 : 16] = ram_temp_output_data[335 : 328];
    compute_data_in_9[31 : 24] = ram_temp_output_data[463 : 456];
    compute_data_in_9[39 : 32] = ram_temp_output_data[591 : 584];
    compute_data_in_9[47 : 40] = ram_temp_output_data[719 : 712];
    compute_data_in_9[55 : 48] = ram_temp_output_data[847 : 840];
    compute_data_in_9[63 : 56] = ram_temp_output_data[975 : 968];
    compute_data_in_9[71 : 64] = ram_temp_output_data[1103 : 1096];
  end

  always @(*) begin
    compute_data_in_10[7 : 0] = ram_temp_output_data[87 : 80];
    compute_data_in_10[15 : 8] = ram_temp_output_data[215 : 208];
    compute_data_in_10[23 : 16] = ram_temp_output_data[343 : 336];
    compute_data_in_10[31 : 24] = ram_temp_output_data[471 : 464];
    compute_data_in_10[39 : 32] = ram_temp_output_data[599 : 592];
    compute_data_in_10[47 : 40] = ram_temp_output_data[727 : 720];
    compute_data_in_10[55 : 48] = ram_temp_output_data[855 : 848];
    compute_data_in_10[63 : 56] = ram_temp_output_data[983 : 976];
    compute_data_in_10[71 : 64] = ram_temp_output_data[1111 : 1104];
  end

  always @(*) begin
    compute_data_in_11[7 : 0] = ram_temp_output_data[95 : 88];
    compute_data_in_11[15 : 8] = ram_temp_output_data[223 : 216];
    compute_data_in_11[23 : 16] = ram_temp_output_data[351 : 344];
    compute_data_in_11[31 : 24] = ram_temp_output_data[479 : 472];
    compute_data_in_11[39 : 32] = ram_temp_output_data[607 : 600];
    compute_data_in_11[47 : 40] = ram_temp_output_data[735 : 728];
    compute_data_in_11[55 : 48] = ram_temp_output_data[863 : 856];
    compute_data_in_11[63 : 56] = ram_temp_output_data[991 : 984];
    compute_data_in_11[71 : 64] = ram_temp_output_data[1119 : 1112];
  end

  always @(*) begin
    compute_data_in_12[7 : 0] = ram_temp_output_data[103 : 96];
    compute_data_in_12[15 : 8] = ram_temp_output_data[231 : 224];
    compute_data_in_12[23 : 16] = ram_temp_output_data[359 : 352];
    compute_data_in_12[31 : 24] = ram_temp_output_data[487 : 480];
    compute_data_in_12[39 : 32] = ram_temp_output_data[615 : 608];
    compute_data_in_12[47 : 40] = ram_temp_output_data[743 : 736];
    compute_data_in_12[55 : 48] = ram_temp_output_data[871 : 864];
    compute_data_in_12[63 : 56] = ram_temp_output_data[999 : 992];
    compute_data_in_12[71 : 64] = ram_temp_output_data[1127 : 1120];
  end

  always @(*) begin
    compute_data_in_13[7 : 0] = ram_temp_output_data[111 : 104];
    compute_data_in_13[15 : 8] = ram_temp_output_data[239 : 232];
    compute_data_in_13[23 : 16] = ram_temp_output_data[367 : 360];
    compute_data_in_13[31 : 24] = ram_temp_output_data[495 : 488];
    compute_data_in_13[39 : 32] = ram_temp_output_data[623 : 616];
    compute_data_in_13[47 : 40] = ram_temp_output_data[751 : 744];
    compute_data_in_13[55 : 48] = ram_temp_output_data[879 : 872];
    compute_data_in_13[63 : 56] = ram_temp_output_data[1007 : 1000];
    compute_data_in_13[71 : 64] = ram_temp_output_data[1135 : 1128];
  end

  always @(*) begin
    compute_data_in_14[7 : 0] = ram_temp_output_data[119 : 112];
    compute_data_in_14[15 : 8] = ram_temp_output_data[247 : 240];
    compute_data_in_14[23 : 16] = ram_temp_output_data[375 : 368];
    compute_data_in_14[31 : 24] = ram_temp_output_data[503 : 496];
    compute_data_in_14[39 : 32] = ram_temp_output_data[631 : 624];
    compute_data_in_14[47 : 40] = ram_temp_output_data[759 : 752];
    compute_data_in_14[55 : 48] = ram_temp_output_data[887 : 880];
    compute_data_in_14[63 : 56] = ram_temp_output_data[1015 : 1008];
    compute_data_in_14[71 : 64] = ram_temp_output_data[1143 : 1136];
  end

  always @(*) begin
    compute_data_in_15[7 : 0] = ram_temp_output_data[127 : 120];
    compute_data_in_15[15 : 8] = ram_temp_output_data[255 : 248];
    compute_data_in_15[23 : 16] = ram_temp_output_data[383 : 376];
    compute_data_in_15[31 : 24] = ram_temp_output_data[511 : 504];
    compute_data_in_15[39 : 32] = ram_temp_output_data[639 : 632];
    compute_data_in_15[47 : 40] = ram_temp_output_data[767 : 760];
    compute_data_in_15[55 : 48] = ram_temp_output_data[895 : 888];
    compute_data_in_15[63 : 56] = ram_temp_output_data[1023 : 1016];
    compute_data_in_15[71 : 64] = ram_temp_output_data[1151 : 1144];
  end

  always @(*) begin
    compute_weight_in_0[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_0[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_0[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_0[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_0[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_0[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_0[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_0[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_0[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_0[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_0[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_0[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_0[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_0[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_0[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_0[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_0[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_0[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_0[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_0[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_0[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_0[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_0[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_0[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_0[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_0[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_0[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_0[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_0[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_0[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_0[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_0[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_0[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_0[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_0[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_0[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_0[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_0[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_0[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_0[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_0[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_0[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_0[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_0[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_0[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_0[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_0[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_0[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_0[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_0[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_0[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_0[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_0[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_0[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_0[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_0[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_0[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_0[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_0[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_0[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_0[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_0[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_0[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_0[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_0[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_0[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_0[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_0[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_0[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_0[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_0[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_0[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_0[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_0[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_0[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_0[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_0[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_0[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_0[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_0[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_0[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_0[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_0[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_0[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_0[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_0[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_0[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_0[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_0[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_0[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_0[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_0[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_0[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_0[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_0[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_0[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_0[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_0[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_0[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_0[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_0[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_0[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_0[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_0[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_0[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_0[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_0[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_0[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_0[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_0[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_0[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_0[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_0[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_0[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_0[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_0[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_0[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_0[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_0[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_0[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_0[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_0[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_0[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_0[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_0[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_0[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_0[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_0[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_0[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_0[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_0[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_0[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_0[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_0[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_0[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_0[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_0[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_0[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_0[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_0[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_0[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_0[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_0[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_0[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_1[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_1[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_1[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_1[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_1[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_1[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_1[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_1[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_1[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_1[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_1[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_1[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_1[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_1[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_1[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_1[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_1[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_1[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_1[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_1[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_1[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_1[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_1[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_1[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_1[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_1[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_1[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_1[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_1[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_1[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_1[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_1[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_1[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_1[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_1[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_1[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_1[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_1[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_1[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_1[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_1[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_1[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_1[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_1[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_1[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_1[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_1[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_1[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_1[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_1[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_1[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_1[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_1[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_1[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_1[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_1[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_1[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_1[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_1[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_1[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_1[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_1[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_1[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_1[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_1[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_1[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_1[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_1[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_1[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_1[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_1[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_1[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_1[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_1[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_1[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_1[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_1[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_1[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_1[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_1[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_1[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_1[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_1[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_1[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_1[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_1[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_1[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_1[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_1[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_1[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_1[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_1[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_1[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_1[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_1[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_1[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_1[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_1[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_1[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_1[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_1[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_1[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_1[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_1[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_1[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_1[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_1[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_1[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_1[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_1[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_1[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_1[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_1[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_1[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_1[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_1[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_1[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_1[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_1[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_1[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_1[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_1[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_1[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_1[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_1[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_1[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_1[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_1[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_1[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_1[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_1[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_1[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_1[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_1[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_1[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_1[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_1[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_1[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_1[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_1[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_1[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_1[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_1[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_1[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_2[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_2[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_2[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_2[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_2[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_2[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_2[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_2[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_2[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_2[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_2[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_2[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_2[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_2[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_2[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_2[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_2[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_2[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_2[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_2[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_2[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_2[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_2[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_2[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_2[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_2[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_2[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_2[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_2[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_2[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_2[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_2[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_2[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_2[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_2[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_2[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_2[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_2[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_2[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_2[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_2[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_2[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_2[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_2[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_2[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_2[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_2[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_2[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_2[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_2[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_2[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_2[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_2[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_2[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_2[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_2[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_2[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_2[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_2[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_2[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_2[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_2[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_2[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_2[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_2[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_2[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_2[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_2[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_2[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_2[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_2[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_2[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_2[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_2[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_2[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_2[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_2[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_2[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_2[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_2[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_2[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_2[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_2[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_2[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_2[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_2[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_2[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_2[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_2[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_2[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_2[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_2[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_2[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_2[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_2[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_2[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_2[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_2[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_2[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_2[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_2[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_2[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_2[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_2[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_2[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_2[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_2[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_2[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_2[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_2[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_2[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_2[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_2[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_2[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_2[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_2[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_2[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_2[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_2[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_2[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_2[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_2[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_2[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_2[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_2[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_2[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_2[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_2[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_2[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_2[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_2[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_2[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_2[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_2[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_2[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_2[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_2[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_2[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_2[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_2[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_2[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_2[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_2[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_2[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_3[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_3[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_3[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_3[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_3[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_3[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_3[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_3[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_3[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_3[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_3[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_3[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_3[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_3[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_3[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_3[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_3[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_3[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_3[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_3[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_3[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_3[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_3[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_3[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_3[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_3[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_3[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_3[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_3[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_3[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_3[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_3[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_3[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_3[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_3[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_3[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_3[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_3[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_3[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_3[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_3[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_3[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_3[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_3[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_3[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_3[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_3[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_3[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_3[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_3[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_3[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_3[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_3[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_3[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_3[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_3[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_3[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_3[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_3[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_3[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_3[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_3[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_3[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_3[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_3[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_3[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_3[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_3[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_3[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_3[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_3[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_3[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_3[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_3[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_3[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_3[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_3[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_3[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_3[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_3[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_3[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_3[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_3[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_3[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_3[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_3[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_3[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_3[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_3[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_3[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_3[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_3[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_3[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_3[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_3[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_3[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_3[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_3[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_3[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_3[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_3[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_3[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_3[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_3[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_3[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_3[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_3[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_3[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_3[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_3[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_3[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_3[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_3[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_3[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_3[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_3[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_3[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_3[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_3[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_3[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_3[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_3[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_3[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_3[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_3[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_3[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_3[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_3[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_3[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_3[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_3[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_3[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_3[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_3[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_3[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_3[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_3[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_3[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_3[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_3[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_3[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_3[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_3[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_3[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_4[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_4[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_4[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_4[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_4[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_4[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_4[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_4[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_4[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_4[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_4[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_4[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_4[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_4[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_4[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_4[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_4[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_4[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_4[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_4[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_4[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_4[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_4[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_4[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_4[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_4[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_4[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_4[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_4[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_4[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_4[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_4[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_4[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_4[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_4[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_4[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_4[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_4[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_4[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_4[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_4[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_4[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_4[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_4[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_4[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_4[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_4[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_4[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_4[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_4[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_4[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_4[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_4[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_4[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_4[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_4[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_4[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_4[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_4[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_4[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_4[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_4[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_4[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_4[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_4[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_4[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_4[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_4[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_4[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_4[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_4[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_4[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_4[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_4[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_4[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_4[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_4[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_4[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_4[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_4[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_4[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_4[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_4[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_4[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_4[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_4[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_4[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_4[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_4[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_4[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_4[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_4[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_4[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_4[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_4[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_4[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_4[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_4[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_4[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_4[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_4[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_4[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_4[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_4[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_4[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_4[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_4[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_4[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_4[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_4[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_4[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_4[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_4[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_4[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_4[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_4[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_4[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_4[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_4[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_4[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_4[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_4[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_4[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_4[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_4[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_4[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_4[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_4[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_4[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_4[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_4[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_4[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_4[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_4[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_4[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_4[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_4[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_4[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_4[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_4[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_4[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_4[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_4[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_4[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_5[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_5[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_5[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_5[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_5[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_5[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_5[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_5[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_5[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_5[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_5[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_5[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_5[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_5[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_5[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_5[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_5[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_5[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_5[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_5[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_5[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_5[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_5[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_5[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_5[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_5[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_5[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_5[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_5[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_5[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_5[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_5[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_5[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_5[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_5[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_5[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_5[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_5[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_5[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_5[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_5[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_5[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_5[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_5[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_5[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_5[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_5[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_5[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_5[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_5[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_5[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_5[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_5[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_5[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_5[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_5[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_5[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_5[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_5[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_5[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_5[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_5[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_5[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_5[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_5[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_5[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_5[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_5[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_5[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_5[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_5[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_5[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_5[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_5[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_5[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_5[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_5[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_5[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_5[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_5[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_5[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_5[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_5[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_5[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_5[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_5[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_5[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_5[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_5[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_5[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_5[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_5[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_5[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_5[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_5[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_5[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_5[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_5[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_5[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_5[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_5[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_5[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_5[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_5[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_5[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_5[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_5[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_5[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_5[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_5[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_5[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_5[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_5[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_5[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_5[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_5[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_5[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_5[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_5[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_5[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_5[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_5[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_5[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_5[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_5[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_5[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_5[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_5[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_5[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_5[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_5[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_5[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_5[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_5[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_5[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_5[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_5[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_5[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_5[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_5[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_5[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_5[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_5[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_5[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_6[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_6[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_6[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_6[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_6[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_6[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_6[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_6[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_6[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_6[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_6[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_6[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_6[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_6[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_6[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_6[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_6[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_6[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_6[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_6[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_6[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_6[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_6[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_6[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_6[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_6[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_6[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_6[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_6[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_6[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_6[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_6[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_6[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_6[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_6[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_6[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_6[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_6[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_6[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_6[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_6[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_6[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_6[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_6[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_6[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_6[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_6[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_6[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_6[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_6[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_6[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_6[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_6[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_6[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_6[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_6[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_6[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_6[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_6[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_6[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_6[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_6[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_6[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_6[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_6[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_6[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_6[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_6[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_6[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_6[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_6[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_6[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_6[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_6[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_6[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_6[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_6[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_6[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_6[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_6[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_6[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_6[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_6[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_6[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_6[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_6[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_6[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_6[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_6[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_6[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_6[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_6[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_6[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_6[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_6[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_6[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_6[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_6[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_6[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_6[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_6[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_6[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_6[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_6[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_6[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_6[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_6[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_6[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_6[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_6[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_6[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_6[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_6[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_6[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_6[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_6[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_6[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_6[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_6[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_6[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_6[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_6[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_6[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_6[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_6[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_6[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_6[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_6[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_6[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_6[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_6[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_6[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_6[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_6[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_6[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_6[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_6[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_6[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_6[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_6[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_6[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_6[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_6[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_6[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  always @(*) begin
    compute_weight_in_7[7 : 0] = load_weight_1_Data_Out_Weight_0[7 : 0];
    compute_weight_in_7[15 : 8] = load_weight_1_Data_Out_Weight_1[7 : 0];
    compute_weight_in_7[23 : 16] = load_weight_1_Data_Out_Weight_2[7 : 0];
    compute_weight_in_7[31 : 24] = load_weight_1_Data_Out_Weight_3[7 : 0];
    compute_weight_in_7[39 : 32] = load_weight_1_Data_Out_Weight_4[7 : 0];
    compute_weight_in_7[47 : 40] = load_weight_1_Data_Out_Weight_5[7 : 0];
    compute_weight_in_7[55 : 48] = load_weight_1_Data_Out_Weight_6[7 : 0];
    compute_weight_in_7[63 : 56] = load_weight_1_Data_Out_Weight_7[7 : 0];
    compute_weight_in_7[71 : 64] = load_weight_1_Data_Out_Weight_8[7 : 0];
    compute_weight_in_7[79 : 72] = load_weight_1_Data_Out_Weight_0[15 : 8];
    compute_weight_in_7[87 : 80] = load_weight_1_Data_Out_Weight_1[15 : 8];
    compute_weight_in_7[95 : 88] = load_weight_1_Data_Out_Weight_2[15 : 8];
    compute_weight_in_7[103 : 96] = load_weight_1_Data_Out_Weight_3[15 : 8];
    compute_weight_in_7[111 : 104] = load_weight_1_Data_Out_Weight_4[15 : 8];
    compute_weight_in_7[119 : 112] = load_weight_1_Data_Out_Weight_5[15 : 8];
    compute_weight_in_7[127 : 120] = load_weight_1_Data_Out_Weight_6[15 : 8];
    compute_weight_in_7[135 : 128] = load_weight_1_Data_Out_Weight_7[15 : 8];
    compute_weight_in_7[143 : 136] = load_weight_1_Data_Out_Weight_8[15 : 8];
    compute_weight_in_7[151 : 144] = load_weight_1_Data_Out_Weight_0[23 : 16];
    compute_weight_in_7[159 : 152] = load_weight_1_Data_Out_Weight_1[23 : 16];
    compute_weight_in_7[167 : 160] = load_weight_1_Data_Out_Weight_2[23 : 16];
    compute_weight_in_7[175 : 168] = load_weight_1_Data_Out_Weight_3[23 : 16];
    compute_weight_in_7[183 : 176] = load_weight_1_Data_Out_Weight_4[23 : 16];
    compute_weight_in_7[191 : 184] = load_weight_1_Data_Out_Weight_5[23 : 16];
    compute_weight_in_7[199 : 192] = load_weight_1_Data_Out_Weight_6[23 : 16];
    compute_weight_in_7[207 : 200] = load_weight_1_Data_Out_Weight_7[23 : 16];
    compute_weight_in_7[215 : 208] = load_weight_1_Data_Out_Weight_8[23 : 16];
    compute_weight_in_7[223 : 216] = load_weight_1_Data_Out_Weight_0[31 : 24];
    compute_weight_in_7[231 : 224] = load_weight_1_Data_Out_Weight_1[31 : 24];
    compute_weight_in_7[239 : 232] = load_weight_1_Data_Out_Weight_2[31 : 24];
    compute_weight_in_7[247 : 240] = load_weight_1_Data_Out_Weight_3[31 : 24];
    compute_weight_in_7[255 : 248] = load_weight_1_Data_Out_Weight_4[31 : 24];
    compute_weight_in_7[263 : 256] = load_weight_1_Data_Out_Weight_5[31 : 24];
    compute_weight_in_7[271 : 264] = load_weight_1_Data_Out_Weight_6[31 : 24];
    compute_weight_in_7[279 : 272] = load_weight_1_Data_Out_Weight_7[31 : 24];
    compute_weight_in_7[287 : 280] = load_weight_1_Data_Out_Weight_8[31 : 24];
    compute_weight_in_7[295 : 288] = load_weight_1_Data_Out_Weight_0[39 : 32];
    compute_weight_in_7[303 : 296] = load_weight_1_Data_Out_Weight_1[39 : 32];
    compute_weight_in_7[311 : 304] = load_weight_1_Data_Out_Weight_2[39 : 32];
    compute_weight_in_7[319 : 312] = load_weight_1_Data_Out_Weight_3[39 : 32];
    compute_weight_in_7[327 : 320] = load_weight_1_Data_Out_Weight_4[39 : 32];
    compute_weight_in_7[335 : 328] = load_weight_1_Data_Out_Weight_5[39 : 32];
    compute_weight_in_7[343 : 336] = load_weight_1_Data_Out_Weight_6[39 : 32];
    compute_weight_in_7[351 : 344] = load_weight_1_Data_Out_Weight_7[39 : 32];
    compute_weight_in_7[359 : 352] = load_weight_1_Data_Out_Weight_8[39 : 32];
    compute_weight_in_7[367 : 360] = load_weight_1_Data_Out_Weight_0[47 : 40];
    compute_weight_in_7[375 : 368] = load_weight_1_Data_Out_Weight_1[47 : 40];
    compute_weight_in_7[383 : 376] = load_weight_1_Data_Out_Weight_2[47 : 40];
    compute_weight_in_7[391 : 384] = load_weight_1_Data_Out_Weight_3[47 : 40];
    compute_weight_in_7[399 : 392] = load_weight_1_Data_Out_Weight_4[47 : 40];
    compute_weight_in_7[407 : 400] = load_weight_1_Data_Out_Weight_5[47 : 40];
    compute_weight_in_7[415 : 408] = load_weight_1_Data_Out_Weight_6[47 : 40];
    compute_weight_in_7[423 : 416] = load_weight_1_Data_Out_Weight_7[47 : 40];
    compute_weight_in_7[431 : 424] = load_weight_1_Data_Out_Weight_8[47 : 40];
    compute_weight_in_7[439 : 432] = load_weight_1_Data_Out_Weight_0[55 : 48];
    compute_weight_in_7[447 : 440] = load_weight_1_Data_Out_Weight_1[55 : 48];
    compute_weight_in_7[455 : 448] = load_weight_1_Data_Out_Weight_2[55 : 48];
    compute_weight_in_7[463 : 456] = load_weight_1_Data_Out_Weight_3[55 : 48];
    compute_weight_in_7[471 : 464] = load_weight_1_Data_Out_Weight_4[55 : 48];
    compute_weight_in_7[479 : 472] = load_weight_1_Data_Out_Weight_5[55 : 48];
    compute_weight_in_7[487 : 480] = load_weight_1_Data_Out_Weight_6[55 : 48];
    compute_weight_in_7[495 : 488] = load_weight_1_Data_Out_Weight_7[55 : 48];
    compute_weight_in_7[503 : 496] = load_weight_1_Data_Out_Weight_8[55 : 48];
    compute_weight_in_7[511 : 504] = load_weight_1_Data_Out_Weight_0[63 : 56];
    compute_weight_in_7[519 : 512] = load_weight_1_Data_Out_Weight_1[63 : 56];
    compute_weight_in_7[527 : 520] = load_weight_1_Data_Out_Weight_2[63 : 56];
    compute_weight_in_7[535 : 528] = load_weight_1_Data_Out_Weight_3[63 : 56];
    compute_weight_in_7[543 : 536] = load_weight_1_Data_Out_Weight_4[63 : 56];
    compute_weight_in_7[551 : 544] = load_weight_1_Data_Out_Weight_5[63 : 56];
    compute_weight_in_7[559 : 552] = load_weight_1_Data_Out_Weight_6[63 : 56];
    compute_weight_in_7[567 : 560] = load_weight_1_Data_Out_Weight_7[63 : 56];
    compute_weight_in_7[575 : 568] = load_weight_1_Data_Out_Weight_8[63 : 56];
    compute_weight_in_7[583 : 576] = load_weight_1_Data_Out_Weight_0[71 : 64];
    compute_weight_in_7[591 : 584] = load_weight_1_Data_Out_Weight_1[71 : 64];
    compute_weight_in_7[599 : 592] = load_weight_1_Data_Out_Weight_2[71 : 64];
    compute_weight_in_7[607 : 600] = load_weight_1_Data_Out_Weight_3[71 : 64];
    compute_weight_in_7[615 : 608] = load_weight_1_Data_Out_Weight_4[71 : 64];
    compute_weight_in_7[623 : 616] = load_weight_1_Data_Out_Weight_5[71 : 64];
    compute_weight_in_7[631 : 624] = load_weight_1_Data_Out_Weight_6[71 : 64];
    compute_weight_in_7[639 : 632] = load_weight_1_Data_Out_Weight_7[71 : 64];
    compute_weight_in_7[647 : 640] = load_weight_1_Data_Out_Weight_8[71 : 64];
    compute_weight_in_7[655 : 648] = load_weight_1_Data_Out_Weight_0[79 : 72];
    compute_weight_in_7[663 : 656] = load_weight_1_Data_Out_Weight_1[79 : 72];
    compute_weight_in_7[671 : 664] = load_weight_1_Data_Out_Weight_2[79 : 72];
    compute_weight_in_7[679 : 672] = load_weight_1_Data_Out_Weight_3[79 : 72];
    compute_weight_in_7[687 : 680] = load_weight_1_Data_Out_Weight_4[79 : 72];
    compute_weight_in_7[695 : 688] = load_weight_1_Data_Out_Weight_5[79 : 72];
    compute_weight_in_7[703 : 696] = load_weight_1_Data_Out_Weight_6[79 : 72];
    compute_weight_in_7[711 : 704] = load_weight_1_Data_Out_Weight_7[79 : 72];
    compute_weight_in_7[719 : 712] = load_weight_1_Data_Out_Weight_8[79 : 72];
    compute_weight_in_7[727 : 720] = load_weight_1_Data_Out_Weight_0[87 : 80];
    compute_weight_in_7[735 : 728] = load_weight_1_Data_Out_Weight_1[87 : 80];
    compute_weight_in_7[743 : 736] = load_weight_1_Data_Out_Weight_2[87 : 80];
    compute_weight_in_7[751 : 744] = load_weight_1_Data_Out_Weight_3[87 : 80];
    compute_weight_in_7[759 : 752] = load_weight_1_Data_Out_Weight_4[87 : 80];
    compute_weight_in_7[767 : 760] = load_weight_1_Data_Out_Weight_5[87 : 80];
    compute_weight_in_7[775 : 768] = load_weight_1_Data_Out_Weight_6[87 : 80];
    compute_weight_in_7[783 : 776] = load_weight_1_Data_Out_Weight_7[87 : 80];
    compute_weight_in_7[791 : 784] = load_weight_1_Data_Out_Weight_8[87 : 80];
    compute_weight_in_7[799 : 792] = load_weight_1_Data_Out_Weight_0[95 : 88];
    compute_weight_in_7[807 : 800] = load_weight_1_Data_Out_Weight_1[95 : 88];
    compute_weight_in_7[815 : 808] = load_weight_1_Data_Out_Weight_2[95 : 88];
    compute_weight_in_7[823 : 816] = load_weight_1_Data_Out_Weight_3[95 : 88];
    compute_weight_in_7[831 : 824] = load_weight_1_Data_Out_Weight_4[95 : 88];
    compute_weight_in_7[839 : 832] = load_weight_1_Data_Out_Weight_5[95 : 88];
    compute_weight_in_7[847 : 840] = load_weight_1_Data_Out_Weight_6[95 : 88];
    compute_weight_in_7[855 : 848] = load_weight_1_Data_Out_Weight_7[95 : 88];
    compute_weight_in_7[863 : 856] = load_weight_1_Data_Out_Weight_8[95 : 88];
    compute_weight_in_7[871 : 864] = load_weight_1_Data_Out_Weight_0[103 : 96];
    compute_weight_in_7[879 : 872] = load_weight_1_Data_Out_Weight_1[103 : 96];
    compute_weight_in_7[887 : 880] = load_weight_1_Data_Out_Weight_2[103 : 96];
    compute_weight_in_7[895 : 888] = load_weight_1_Data_Out_Weight_3[103 : 96];
    compute_weight_in_7[903 : 896] = load_weight_1_Data_Out_Weight_4[103 : 96];
    compute_weight_in_7[911 : 904] = load_weight_1_Data_Out_Weight_5[103 : 96];
    compute_weight_in_7[919 : 912] = load_weight_1_Data_Out_Weight_6[103 : 96];
    compute_weight_in_7[927 : 920] = load_weight_1_Data_Out_Weight_7[103 : 96];
    compute_weight_in_7[935 : 928] = load_weight_1_Data_Out_Weight_8[103 : 96];
    compute_weight_in_7[943 : 936] = load_weight_1_Data_Out_Weight_0[111 : 104];
    compute_weight_in_7[951 : 944] = load_weight_1_Data_Out_Weight_1[111 : 104];
    compute_weight_in_7[959 : 952] = load_weight_1_Data_Out_Weight_2[111 : 104];
    compute_weight_in_7[967 : 960] = load_weight_1_Data_Out_Weight_3[111 : 104];
    compute_weight_in_7[975 : 968] = load_weight_1_Data_Out_Weight_4[111 : 104];
    compute_weight_in_7[983 : 976] = load_weight_1_Data_Out_Weight_5[111 : 104];
    compute_weight_in_7[991 : 984] = load_weight_1_Data_Out_Weight_6[111 : 104];
    compute_weight_in_7[999 : 992] = load_weight_1_Data_Out_Weight_7[111 : 104];
    compute_weight_in_7[1007 : 1000] = load_weight_1_Data_Out_Weight_8[111 : 104];
    compute_weight_in_7[1015 : 1008] = load_weight_1_Data_Out_Weight_0[119 : 112];
    compute_weight_in_7[1023 : 1016] = load_weight_1_Data_Out_Weight_1[119 : 112];
    compute_weight_in_7[1031 : 1024] = load_weight_1_Data_Out_Weight_2[119 : 112];
    compute_weight_in_7[1039 : 1032] = load_weight_1_Data_Out_Weight_3[119 : 112];
    compute_weight_in_7[1047 : 1040] = load_weight_1_Data_Out_Weight_4[119 : 112];
    compute_weight_in_7[1055 : 1048] = load_weight_1_Data_Out_Weight_5[119 : 112];
    compute_weight_in_7[1063 : 1056] = load_weight_1_Data_Out_Weight_6[119 : 112];
    compute_weight_in_7[1071 : 1064] = load_weight_1_Data_Out_Weight_7[119 : 112];
    compute_weight_in_7[1079 : 1072] = load_weight_1_Data_Out_Weight_8[119 : 112];
    compute_weight_in_7[1087 : 1080] = load_weight_1_Data_Out_Weight_0[127 : 120];
    compute_weight_in_7[1095 : 1088] = load_weight_1_Data_Out_Weight_1[127 : 120];
    compute_weight_in_7[1103 : 1096] = load_weight_1_Data_Out_Weight_2[127 : 120];
    compute_weight_in_7[1111 : 1104] = load_weight_1_Data_Out_Weight_3[127 : 120];
    compute_weight_in_7[1119 : 1112] = load_weight_1_Data_Out_Weight_4[127 : 120];
    compute_weight_in_7[1127 : 1120] = load_weight_1_Data_Out_Weight_5[127 : 120];
    compute_weight_in_7[1135 : 1128] = load_weight_1_Data_Out_Weight_6[127 : 120];
    compute_weight_in_7[1143 : 1136] = load_weight_1_Data_Out_Weight_7[127 : 120];
    compute_weight_in_7[1151 : 1144] = load_weight_1_Data_Out_Weight_8[127 : 120];
  end

  assign compute_weight_in_delay_0 = compute_weight_in_0_regNext;
  assign compute_weight_in_delay_1 = compute_weight_in_1_regNext;
  assign compute_weight_in_delay_2 = compute_weight_in_2_regNext;
  assign compute_weight_in_delay_3 = compute_weight_in_3_regNext;
  assign compute_weight_in_delay_4 = compute_weight_in_4_regNext;
  assign compute_weight_in_delay_5 = compute_weight_in_5_regNext;
  assign compute_weight_in_delay_6 = compute_weight_in_6_regNext;
  assign compute_weight_in_delay_7 = compute_weight_in_7_regNext;
  assign mul_add_simd_128_weightIn = compute_weight_in_0[71 : 0];
  always @(*) begin
    compute_data_out_0[19 : 0] = mul_add_simd_128_dataOut;
    compute_data_out_0[39 : 20] = mul_add_simd_129_dataOut;
    compute_data_out_0[59 : 40] = mul_add_simd_130_dataOut;
    compute_data_out_0[79 : 60] = mul_add_simd_131_dataOut;
    compute_data_out_0[99 : 80] = mul_add_simd_132_dataOut;
    compute_data_out_0[119 : 100] = mul_add_simd_133_dataOut;
    compute_data_out_0[139 : 120] = mul_add_simd_134_dataOut;
    compute_data_out_0[159 : 140] = mul_add_simd_135_dataOut;
    compute_data_out_0[179 : 160] = mul_add_simd_136_dataOut;
    compute_data_out_0[199 : 180] = mul_add_simd_137_dataOut;
    compute_data_out_0[219 : 200] = mul_add_simd_138_dataOut;
    compute_data_out_0[239 : 220] = mul_add_simd_139_dataOut;
    compute_data_out_0[259 : 240] = mul_add_simd_140_dataOut;
    compute_data_out_0[279 : 260] = mul_add_simd_141_dataOut;
    compute_data_out_0[299 : 280] = mul_add_simd_142_dataOut;
    compute_data_out_0[319 : 300] = mul_add_simd_143_dataOut;
  end

  assign mul_add_simd_129_weightIn = compute_weight_in_0[143 : 72];
  assign mul_add_simd_130_weightIn = compute_weight_in_0[215 : 144];
  assign mul_add_simd_131_weightIn = compute_weight_in_0[287 : 216];
  assign mul_add_simd_132_weightIn = compute_weight_in_0[359 : 288];
  assign mul_add_simd_133_weightIn = compute_weight_in_0[431 : 360];
  assign mul_add_simd_134_weightIn = compute_weight_in_0[503 : 432];
  assign mul_add_simd_135_weightIn = compute_weight_in_0[575 : 504];
  assign mul_add_simd_136_weightIn = compute_weight_in_0[647 : 576];
  assign mul_add_simd_137_weightIn = compute_weight_in_0[719 : 648];
  assign mul_add_simd_138_weightIn = compute_weight_in_0[791 : 720];
  assign mul_add_simd_139_weightIn = compute_weight_in_0[863 : 792];
  assign mul_add_simd_140_weightIn = compute_weight_in_0[935 : 864];
  assign mul_add_simd_141_weightIn = compute_weight_in_0[1007 : 936];
  assign mul_add_simd_142_weightIn = compute_weight_in_0[1079 : 1008];
  assign mul_add_simd_143_weightIn = compute_weight_in_0[1151 : 1080];
  assign mul_add_simd_144_weightIn = compute_weight_in_1[71 : 0];
  always @(*) begin
    compute_data_out_1[19 : 0] = mul_add_simd_144_dataOut;
    compute_data_out_1[39 : 20] = mul_add_simd_145_dataOut;
    compute_data_out_1[59 : 40] = mul_add_simd_146_dataOut;
    compute_data_out_1[79 : 60] = mul_add_simd_147_dataOut;
    compute_data_out_1[99 : 80] = mul_add_simd_148_dataOut;
    compute_data_out_1[119 : 100] = mul_add_simd_149_dataOut;
    compute_data_out_1[139 : 120] = mul_add_simd_150_dataOut;
    compute_data_out_1[159 : 140] = mul_add_simd_151_dataOut;
    compute_data_out_1[179 : 160] = mul_add_simd_152_dataOut;
    compute_data_out_1[199 : 180] = mul_add_simd_153_dataOut;
    compute_data_out_1[219 : 200] = mul_add_simd_154_dataOut;
    compute_data_out_1[239 : 220] = mul_add_simd_155_dataOut;
    compute_data_out_1[259 : 240] = mul_add_simd_156_dataOut;
    compute_data_out_1[279 : 260] = mul_add_simd_157_dataOut;
    compute_data_out_1[299 : 280] = mul_add_simd_158_dataOut;
    compute_data_out_1[319 : 300] = mul_add_simd_159_dataOut;
  end

  assign mul_add_simd_145_weightIn = compute_weight_in_1[143 : 72];
  assign mul_add_simd_146_weightIn = compute_weight_in_1[215 : 144];
  assign mul_add_simd_147_weightIn = compute_weight_in_1[287 : 216];
  assign mul_add_simd_148_weightIn = compute_weight_in_1[359 : 288];
  assign mul_add_simd_149_weightIn = compute_weight_in_1[431 : 360];
  assign mul_add_simd_150_weightIn = compute_weight_in_1[503 : 432];
  assign mul_add_simd_151_weightIn = compute_weight_in_1[575 : 504];
  assign mul_add_simd_152_weightIn = compute_weight_in_1[647 : 576];
  assign mul_add_simd_153_weightIn = compute_weight_in_1[719 : 648];
  assign mul_add_simd_154_weightIn = compute_weight_in_1[791 : 720];
  assign mul_add_simd_155_weightIn = compute_weight_in_1[863 : 792];
  assign mul_add_simd_156_weightIn = compute_weight_in_1[935 : 864];
  assign mul_add_simd_157_weightIn = compute_weight_in_1[1007 : 936];
  assign mul_add_simd_158_weightIn = compute_weight_in_1[1079 : 1008];
  assign mul_add_simd_159_weightIn = compute_weight_in_1[1151 : 1080];
  assign mul_add_simd_160_weightIn = compute_weight_in_2[71 : 0];
  always @(*) begin
    compute_data_out_2[19 : 0] = mul_add_simd_160_dataOut;
    compute_data_out_2[39 : 20] = mul_add_simd_161_dataOut;
    compute_data_out_2[59 : 40] = mul_add_simd_162_dataOut;
    compute_data_out_2[79 : 60] = mul_add_simd_163_dataOut;
    compute_data_out_2[99 : 80] = mul_add_simd_164_dataOut;
    compute_data_out_2[119 : 100] = mul_add_simd_165_dataOut;
    compute_data_out_2[139 : 120] = mul_add_simd_166_dataOut;
    compute_data_out_2[159 : 140] = mul_add_simd_167_dataOut;
    compute_data_out_2[179 : 160] = mul_add_simd_168_dataOut;
    compute_data_out_2[199 : 180] = mul_add_simd_169_dataOut;
    compute_data_out_2[219 : 200] = mul_add_simd_170_dataOut;
    compute_data_out_2[239 : 220] = mul_add_simd_171_dataOut;
    compute_data_out_2[259 : 240] = mul_add_simd_172_dataOut;
    compute_data_out_2[279 : 260] = mul_add_simd_173_dataOut;
    compute_data_out_2[299 : 280] = mul_add_simd_174_dataOut;
    compute_data_out_2[319 : 300] = mul_add_simd_175_dataOut;
  end

  assign mul_add_simd_161_weightIn = compute_weight_in_2[143 : 72];
  assign mul_add_simd_162_weightIn = compute_weight_in_2[215 : 144];
  assign mul_add_simd_163_weightIn = compute_weight_in_2[287 : 216];
  assign mul_add_simd_164_weightIn = compute_weight_in_2[359 : 288];
  assign mul_add_simd_165_weightIn = compute_weight_in_2[431 : 360];
  assign mul_add_simd_166_weightIn = compute_weight_in_2[503 : 432];
  assign mul_add_simd_167_weightIn = compute_weight_in_2[575 : 504];
  assign mul_add_simd_168_weightIn = compute_weight_in_2[647 : 576];
  assign mul_add_simd_169_weightIn = compute_weight_in_2[719 : 648];
  assign mul_add_simd_170_weightIn = compute_weight_in_2[791 : 720];
  assign mul_add_simd_171_weightIn = compute_weight_in_2[863 : 792];
  assign mul_add_simd_172_weightIn = compute_weight_in_2[935 : 864];
  assign mul_add_simd_173_weightIn = compute_weight_in_2[1007 : 936];
  assign mul_add_simd_174_weightIn = compute_weight_in_2[1079 : 1008];
  assign mul_add_simd_175_weightIn = compute_weight_in_2[1151 : 1080];
  assign mul_add_simd_176_weightIn = compute_weight_in_3[71 : 0];
  always @(*) begin
    compute_data_out_3[19 : 0] = mul_add_simd_176_dataOut;
    compute_data_out_3[39 : 20] = mul_add_simd_177_dataOut;
    compute_data_out_3[59 : 40] = mul_add_simd_178_dataOut;
    compute_data_out_3[79 : 60] = mul_add_simd_179_dataOut;
    compute_data_out_3[99 : 80] = mul_add_simd_180_dataOut;
    compute_data_out_3[119 : 100] = mul_add_simd_181_dataOut;
    compute_data_out_3[139 : 120] = mul_add_simd_182_dataOut;
    compute_data_out_3[159 : 140] = mul_add_simd_183_dataOut;
    compute_data_out_3[179 : 160] = mul_add_simd_184_dataOut;
    compute_data_out_3[199 : 180] = mul_add_simd_185_dataOut;
    compute_data_out_3[219 : 200] = mul_add_simd_186_dataOut;
    compute_data_out_3[239 : 220] = mul_add_simd_187_dataOut;
    compute_data_out_3[259 : 240] = mul_add_simd_188_dataOut;
    compute_data_out_3[279 : 260] = mul_add_simd_189_dataOut;
    compute_data_out_3[299 : 280] = mul_add_simd_190_dataOut;
    compute_data_out_3[319 : 300] = mul_add_simd_191_dataOut;
  end

  assign mul_add_simd_177_weightIn = compute_weight_in_3[143 : 72];
  assign mul_add_simd_178_weightIn = compute_weight_in_3[215 : 144];
  assign mul_add_simd_179_weightIn = compute_weight_in_3[287 : 216];
  assign mul_add_simd_180_weightIn = compute_weight_in_3[359 : 288];
  assign mul_add_simd_181_weightIn = compute_weight_in_3[431 : 360];
  assign mul_add_simd_182_weightIn = compute_weight_in_3[503 : 432];
  assign mul_add_simd_183_weightIn = compute_weight_in_3[575 : 504];
  assign mul_add_simd_184_weightIn = compute_weight_in_3[647 : 576];
  assign mul_add_simd_185_weightIn = compute_weight_in_3[719 : 648];
  assign mul_add_simd_186_weightIn = compute_weight_in_3[791 : 720];
  assign mul_add_simd_187_weightIn = compute_weight_in_3[863 : 792];
  assign mul_add_simd_188_weightIn = compute_weight_in_3[935 : 864];
  assign mul_add_simd_189_weightIn = compute_weight_in_3[1007 : 936];
  assign mul_add_simd_190_weightIn = compute_weight_in_3[1079 : 1008];
  assign mul_add_simd_191_weightIn = compute_weight_in_3[1151 : 1080];
  assign mul_add_simd_192_weightIn = compute_weight_in_4[71 : 0];
  always @(*) begin
    compute_data_out_4[19 : 0] = mul_add_simd_192_dataOut;
    compute_data_out_4[39 : 20] = mul_add_simd_193_dataOut;
    compute_data_out_4[59 : 40] = mul_add_simd_194_dataOut;
    compute_data_out_4[79 : 60] = mul_add_simd_195_dataOut;
    compute_data_out_4[99 : 80] = mul_add_simd_196_dataOut;
    compute_data_out_4[119 : 100] = mul_add_simd_197_dataOut;
    compute_data_out_4[139 : 120] = mul_add_simd_198_dataOut;
    compute_data_out_4[159 : 140] = mul_add_simd_199_dataOut;
    compute_data_out_4[179 : 160] = mul_add_simd_200_dataOut;
    compute_data_out_4[199 : 180] = mul_add_simd_201_dataOut;
    compute_data_out_4[219 : 200] = mul_add_simd_202_dataOut;
    compute_data_out_4[239 : 220] = mul_add_simd_203_dataOut;
    compute_data_out_4[259 : 240] = mul_add_simd_204_dataOut;
    compute_data_out_4[279 : 260] = mul_add_simd_205_dataOut;
    compute_data_out_4[299 : 280] = mul_add_simd_206_dataOut;
    compute_data_out_4[319 : 300] = mul_add_simd_207_dataOut;
  end

  assign mul_add_simd_193_weightIn = compute_weight_in_4[143 : 72];
  assign mul_add_simd_194_weightIn = compute_weight_in_4[215 : 144];
  assign mul_add_simd_195_weightIn = compute_weight_in_4[287 : 216];
  assign mul_add_simd_196_weightIn = compute_weight_in_4[359 : 288];
  assign mul_add_simd_197_weightIn = compute_weight_in_4[431 : 360];
  assign mul_add_simd_198_weightIn = compute_weight_in_4[503 : 432];
  assign mul_add_simd_199_weightIn = compute_weight_in_4[575 : 504];
  assign mul_add_simd_200_weightIn = compute_weight_in_4[647 : 576];
  assign mul_add_simd_201_weightIn = compute_weight_in_4[719 : 648];
  assign mul_add_simd_202_weightIn = compute_weight_in_4[791 : 720];
  assign mul_add_simd_203_weightIn = compute_weight_in_4[863 : 792];
  assign mul_add_simd_204_weightIn = compute_weight_in_4[935 : 864];
  assign mul_add_simd_205_weightIn = compute_weight_in_4[1007 : 936];
  assign mul_add_simd_206_weightIn = compute_weight_in_4[1079 : 1008];
  assign mul_add_simd_207_weightIn = compute_weight_in_4[1151 : 1080];
  assign mul_add_simd_208_weightIn = compute_weight_in_5[71 : 0];
  always @(*) begin
    compute_data_out_5[19 : 0] = mul_add_simd_208_dataOut;
    compute_data_out_5[39 : 20] = mul_add_simd_209_dataOut;
    compute_data_out_5[59 : 40] = mul_add_simd_210_dataOut;
    compute_data_out_5[79 : 60] = mul_add_simd_211_dataOut;
    compute_data_out_5[99 : 80] = mul_add_simd_212_dataOut;
    compute_data_out_5[119 : 100] = mul_add_simd_213_dataOut;
    compute_data_out_5[139 : 120] = mul_add_simd_214_dataOut;
    compute_data_out_5[159 : 140] = mul_add_simd_215_dataOut;
    compute_data_out_5[179 : 160] = mul_add_simd_216_dataOut;
    compute_data_out_5[199 : 180] = mul_add_simd_217_dataOut;
    compute_data_out_5[219 : 200] = mul_add_simd_218_dataOut;
    compute_data_out_5[239 : 220] = mul_add_simd_219_dataOut;
    compute_data_out_5[259 : 240] = mul_add_simd_220_dataOut;
    compute_data_out_5[279 : 260] = mul_add_simd_221_dataOut;
    compute_data_out_5[299 : 280] = mul_add_simd_222_dataOut;
    compute_data_out_5[319 : 300] = mul_add_simd_223_dataOut;
  end

  assign mul_add_simd_209_weightIn = compute_weight_in_5[143 : 72];
  assign mul_add_simd_210_weightIn = compute_weight_in_5[215 : 144];
  assign mul_add_simd_211_weightIn = compute_weight_in_5[287 : 216];
  assign mul_add_simd_212_weightIn = compute_weight_in_5[359 : 288];
  assign mul_add_simd_213_weightIn = compute_weight_in_5[431 : 360];
  assign mul_add_simd_214_weightIn = compute_weight_in_5[503 : 432];
  assign mul_add_simd_215_weightIn = compute_weight_in_5[575 : 504];
  assign mul_add_simd_216_weightIn = compute_weight_in_5[647 : 576];
  assign mul_add_simd_217_weightIn = compute_weight_in_5[719 : 648];
  assign mul_add_simd_218_weightIn = compute_weight_in_5[791 : 720];
  assign mul_add_simd_219_weightIn = compute_weight_in_5[863 : 792];
  assign mul_add_simd_220_weightIn = compute_weight_in_5[935 : 864];
  assign mul_add_simd_221_weightIn = compute_weight_in_5[1007 : 936];
  assign mul_add_simd_222_weightIn = compute_weight_in_5[1079 : 1008];
  assign mul_add_simd_223_weightIn = compute_weight_in_5[1151 : 1080];
  assign mul_add_simd_224_weightIn = compute_weight_in_6[71 : 0];
  always @(*) begin
    compute_data_out_6[19 : 0] = mul_add_simd_224_dataOut;
    compute_data_out_6[39 : 20] = mul_add_simd_225_dataOut;
    compute_data_out_6[59 : 40] = mul_add_simd_226_dataOut;
    compute_data_out_6[79 : 60] = mul_add_simd_227_dataOut;
    compute_data_out_6[99 : 80] = mul_add_simd_228_dataOut;
    compute_data_out_6[119 : 100] = mul_add_simd_229_dataOut;
    compute_data_out_6[139 : 120] = mul_add_simd_230_dataOut;
    compute_data_out_6[159 : 140] = mul_add_simd_231_dataOut;
    compute_data_out_6[179 : 160] = mul_add_simd_232_dataOut;
    compute_data_out_6[199 : 180] = mul_add_simd_233_dataOut;
    compute_data_out_6[219 : 200] = mul_add_simd_234_dataOut;
    compute_data_out_6[239 : 220] = mul_add_simd_235_dataOut;
    compute_data_out_6[259 : 240] = mul_add_simd_236_dataOut;
    compute_data_out_6[279 : 260] = mul_add_simd_237_dataOut;
    compute_data_out_6[299 : 280] = mul_add_simd_238_dataOut;
    compute_data_out_6[319 : 300] = mul_add_simd_239_dataOut;
  end

  assign mul_add_simd_225_weightIn = compute_weight_in_6[143 : 72];
  assign mul_add_simd_226_weightIn = compute_weight_in_6[215 : 144];
  assign mul_add_simd_227_weightIn = compute_weight_in_6[287 : 216];
  assign mul_add_simd_228_weightIn = compute_weight_in_6[359 : 288];
  assign mul_add_simd_229_weightIn = compute_weight_in_6[431 : 360];
  assign mul_add_simd_230_weightIn = compute_weight_in_6[503 : 432];
  assign mul_add_simd_231_weightIn = compute_weight_in_6[575 : 504];
  assign mul_add_simd_232_weightIn = compute_weight_in_6[647 : 576];
  assign mul_add_simd_233_weightIn = compute_weight_in_6[719 : 648];
  assign mul_add_simd_234_weightIn = compute_weight_in_6[791 : 720];
  assign mul_add_simd_235_weightIn = compute_weight_in_6[863 : 792];
  assign mul_add_simd_236_weightIn = compute_weight_in_6[935 : 864];
  assign mul_add_simd_237_weightIn = compute_weight_in_6[1007 : 936];
  assign mul_add_simd_238_weightIn = compute_weight_in_6[1079 : 1008];
  assign mul_add_simd_239_weightIn = compute_weight_in_6[1151 : 1080];
  assign mul_add_simd_240_weightIn = compute_weight_in_7[71 : 0];
  always @(*) begin
    compute_data_out_7[19 : 0] = mul_add_simd_240_dataOut;
    compute_data_out_7[39 : 20] = mul_add_simd_241_dataOut;
    compute_data_out_7[59 : 40] = mul_add_simd_242_dataOut;
    compute_data_out_7[79 : 60] = mul_add_simd_243_dataOut;
    compute_data_out_7[99 : 80] = mul_add_simd_244_dataOut;
    compute_data_out_7[119 : 100] = mul_add_simd_245_dataOut;
    compute_data_out_7[139 : 120] = mul_add_simd_246_dataOut;
    compute_data_out_7[159 : 140] = mul_add_simd_247_dataOut;
    compute_data_out_7[179 : 160] = mul_add_simd_248_dataOut;
    compute_data_out_7[199 : 180] = mul_add_simd_249_dataOut;
    compute_data_out_7[219 : 200] = mul_add_simd_250_dataOut;
    compute_data_out_7[239 : 220] = mul_add_simd_251_dataOut;
    compute_data_out_7[259 : 240] = mul_add_simd_252_dataOut;
    compute_data_out_7[279 : 260] = mul_add_simd_253_dataOut;
    compute_data_out_7[299 : 280] = mul_add_simd_254_dataOut;
    compute_data_out_7[319 : 300] = mul_add_simd_255_dataOut;
  end

  assign mul_add_simd_241_weightIn = compute_weight_in_7[143 : 72];
  assign mul_add_simd_242_weightIn = compute_weight_in_7[215 : 144];
  assign mul_add_simd_243_weightIn = compute_weight_in_7[287 : 216];
  assign mul_add_simd_244_weightIn = compute_weight_in_7[359 : 288];
  assign mul_add_simd_245_weightIn = compute_weight_in_7[431 : 360];
  assign mul_add_simd_246_weightIn = compute_weight_in_7[503 : 432];
  assign mul_add_simd_247_weightIn = compute_weight_in_7[575 : 504];
  assign mul_add_simd_248_weightIn = compute_weight_in_7[647 : 576];
  assign mul_add_simd_249_weightIn = compute_weight_in_7[719 : 648];
  assign mul_add_simd_250_weightIn = compute_weight_in_7[791 : 720];
  assign mul_add_simd_251_weightIn = compute_weight_in_7[863 : 792];
  assign mul_add_simd_252_weightIn = compute_weight_in_7[935 : 864];
  assign mul_add_simd_253_weightIn = compute_weight_in_7[1007 : 936];
  assign mul_add_simd_254_weightIn = compute_weight_in_7[1079 : 1008];
  assign mul_add_simd_255_weightIn = compute_weight_in_7[1151 : 1080];
  assign data_result_temp_0 = channel_in_acc_8_data_out;
  assign data_result_temp_1 = channel_in_acc_9_data_out;
  assign data_result_temp_2 = channel_in_acc_10_data_out;
  assign data_result_temp_3 = channel_in_acc_11_data_out;
  assign data_result_temp_4 = channel_in_acc_12_data_out;
  assign data_result_temp_5 = channel_in_acc_13_data_out;
  assign data_result_temp_6 = channel_in_acc_14_data_out;
  assign data_result_temp_7 = channel_in_acc_15_data_out;
  always @(*) begin
    M_DATA_payload[31 : 0] = channel_out_acc_8_data_out;
    M_DATA_payload[63 : 32] = channel_out_acc_9_data_out;
    M_DATA_payload[95 : 64] = channel_out_acc_10_data_out;
    M_DATA_payload[127 : 96] = channel_out_acc_11_data_out;
    M_DATA_payload[159 : 128] = channel_out_acc_12_data_out;
    M_DATA_payload[191 : 160] = channel_out_acc_13_data_out;
    M_DATA_payload[223 : 192] = channel_out_acc_14_data_out;
    M_DATA_payload[255 : 224] = channel_out_acc_15_data_out;
  end

  always @(posedge clk) begin
    compute_ctrl_1_M_Valid_regNext <= compute_ctrl_1_M_Valid;
    M_DATA_valid <= compute_ctrl_1_M_Valid_regNext;
    ram_temp_output_data_delay_1 <= ram_temp_output_data;
    ram_temp_output_data_delay <= ram_temp_output_data_delay_1;
    compute_weight_in_0_regNext <= compute_weight_in_0;
    compute_weight_in_1_regNext <= compute_weight_in_1;
    compute_weight_in_2_regNext <= compute_weight_in_2;
    compute_weight_in_3_regNext <= compute_weight_in_3;
    compute_weight_in_4_regNext <= compute_weight_in_4;
    compute_weight_in_5_regNext <= compute_weight_in_5;
    compute_weight_in_6_regNext <= compute_weight_in_6;
    compute_weight_in_7_regNext <= compute_weight_in_7;
  end


endmodule
